magic
tech sky130A
magscale 1 2
timestamp 1640967747
<< locali >>
rect 161305 556223 161339 557345
rect 208961 556699 208995 557345
rect 217793 556971 217827 557345
rect 359565 557243 359599 557413
rect 365637 557039 365671 557413
rect 368489 556903 368523 557413
rect 371525 556835 371559 557413
rect 374469 556767 374503 557413
rect 377413 556631 377447 557413
rect 383761 556563 383795 557413
rect 389189 556495 389223 557413
rect 392133 556427 392167 557413
rect 401149 556359 401183 557413
rect 404185 556291 404219 557413
rect 426173 147747 426207 148325
rect 398205 4811 398239 4845
rect 398055 4777 398239 4811
rect 523601 4641 523785 4675
rect 523601 4607 523635 4641
rect 98561 3247 98595 4097
rect 237297 3859 237331 3961
rect 229661 3825 229937 3859
rect 229661 3655 229695 3825
rect 229787 3757 230029 3791
rect 226349 3621 226625 3655
rect 226349 3587 226383 3621
rect 229235 3485 229477 3519
rect 230765 3451 230799 3825
rect 237297 3825 237481 3859
rect 231869 3519 231903 3825
rect 236101 3451 236135 3621
rect 238769 3383 238803 3621
rect 238861 3315 238895 3893
rect 315221 3723 315255 3961
rect 319913 3859 319947 3961
rect 315129 3519 315163 3689
rect 229661 2975 229695 3009
rect 229661 2941 229845 2975
rect 126103 2873 126253 2907
<< viali >>
rect 359565 557413 359599 557447
rect 161305 557345 161339 557379
rect 208961 557345 208995 557379
rect 217793 557345 217827 557379
rect 359565 557209 359599 557243
rect 365637 557413 365671 557447
rect 365637 557005 365671 557039
rect 368489 557413 368523 557447
rect 217793 556937 217827 556971
rect 368489 556869 368523 556903
rect 371525 557413 371559 557447
rect 371525 556801 371559 556835
rect 374469 557413 374503 557447
rect 374469 556733 374503 556767
rect 377413 557413 377447 557447
rect 208961 556665 208995 556699
rect 377413 556597 377447 556631
rect 383761 557413 383795 557447
rect 383761 556529 383795 556563
rect 389189 557413 389223 557447
rect 389189 556461 389223 556495
rect 392133 557413 392167 557447
rect 392133 556393 392167 556427
rect 401149 557413 401183 557447
rect 401149 556325 401183 556359
rect 404185 557413 404219 557447
rect 404185 556257 404219 556291
rect 161305 556189 161339 556223
rect 426173 148325 426207 148359
rect 426173 147713 426207 147747
rect 398205 4845 398239 4879
rect 398021 4777 398055 4811
rect 523785 4641 523819 4675
rect 523601 4573 523635 4607
rect 98561 4097 98595 4131
rect 237297 3961 237331 3995
rect 315221 3961 315255 3995
rect 238861 3893 238895 3927
rect 229937 3825 229971 3859
rect 230765 3825 230799 3859
rect 229753 3757 229787 3791
rect 230029 3757 230063 3791
rect 226625 3621 226659 3655
rect 229661 3621 229695 3655
rect 226349 3553 226383 3587
rect 229201 3485 229235 3519
rect 229477 3485 229511 3519
rect 231869 3825 231903 3859
rect 237481 3825 237515 3859
rect 231869 3485 231903 3519
rect 236101 3621 236135 3655
rect 230765 3417 230799 3451
rect 236101 3417 236135 3451
rect 238769 3621 238803 3655
rect 238769 3349 238803 3383
rect 319913 3961 319947 3995
rect 319913 3825 319947 3859
rect 315129 3689 315163 3723
rect 315221 3689 315255 3723
rect 315129 3485 315163 3519
rect 238861 3281 238895 3315
rect 98561 3213 98595 3247
rect 229661 3009 229695 3043
rect 229845 2941 229879 2975
rect 126069 2873 126103 2907
rect 126253 2873 126287 2907
<< metal1 >>
rect 154114 700952 154120 701004
rect 154172 700992 154178 701004
rect 317414 700992 317420 701004
rect 154172 700964 317420 700992
rect 154172 700952 154178 700964
rect 317414 700952 317420 700964
rect 317472 700952 317478 701004
rect 137830 700884 137836 700936
rect 137888 700924 137894 700936
rect 314654 700924 314660 700936
rect 137888 700896 314660 700924
rect 137888 700884 137894 700896
rect 314654 700884 314660 700896
rect 314712 700884 314718 700936
rect 271782 700816 271788 700868
rect 271840 700856 271846 700868
rect 462314 700856 462320 700868
rect 271840 700828 462320 700856
rect 271840 700816 271846 700828
rect 462314 700816 462320 700828
rect 462372 700816 462378 700868
rect 274542 700748 274548 700800
rect 274600 700788 274606 700800
rect 478506 700788 478512 700800
rect 274600 700760 478512 700788
rect 274600 700748 274606 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 89162 700680 89168 700732
rect 89220 700720 89226 700732
rect 327074 700720 327080 700732
rect 89220 700692 327080 700720
rect 89220 700680 89226 700692
rect 327074 700680 327080 700692
rect 327132 700680 327138 700732
rect 72970 700612 72976 700664
rect 73028 700652 73034 700664
rect 324314 700652 324320 700664
rect 73028 700624 324320 700652
rect 73028 700612 73034 700624
rect 324314 700612 324320 700624
rect 324372 700612 324378 700664
rect 262122 700544 262128 700596
rect 262180 700584 262186 700596
rect 527174 700584 527180 700596
rect 262180 700556 527180 700584
rect 262180 700544 262186 700556
rect 527174 700544 527180 700556
rect 527232 700544 527238 700596
rect 264882 700476 264888 700528
rect 264940 700516 264946 700528
rect 543458 700516 543464 700528
rect 264940 700488 543464 700516
rect 264940 700476 264946 700488
rect 543458 700476 543464 700488
rect 543516 700476 543522 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 329834 700448 329840 700460
rect 40552 700420 329840 700448
rect 40552 700408 40558 700420
rect 329834 700408 329840 700420
rect 329892 700408 329898 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 335354 700380 335360 700392
rect 24360 700352 335360 700380
rect 24360 700340 24366 700352
rect 335354 700340 335360 700352
rect 335412 700340 335418 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 332594 700312 332600 700324
rect 8168 700284 332600 700312
rect 8168 700272 8174 700284
rect 332594 700272 332600 700284
rect 332652 700272 332658 700324
rect 282822 700204 282828 700256
rect 282880 700244 282886 700256
rect 413646 700244 413652 700256
rect 282880 700216 413652 700244
rect 282880 700204 282886 700216
rect 413646 700204 413652 700216
rect 413704 700204 413710 700256
rect 280062 700136 280068 700188
rect 280120 700176 280126 700188
rect 397454 700176 397460 700188
rect 280120 700148 397460 700176
rect 280120 700136 280126 700148
rect 397454 700136 397460 700148
rect 397512 700136 397518 700188
rect 202782 700068 202788 700120
rect 202840 700108 202846 700120
rect 306374 700108 306380 700120
rect 202840 700080 306380 700108
rect 202840 700068 202846 700080
rect 306374 700068 306380 700080
rect 306432 700068 306438 700120
rect 218974 700000 218980 700052
rect 219032 700040 219038 700052
rect 309134 700040 309140 700052
rect 219032 700012 309140 700040
rect 219032 700000 219038 700012
rect 309134 700000 309140 700012
rect 309192 700000 309198 700052
rect 292482 699932 292488 699984
rect 292540 699972 292546 699984
rect 348786 699972 348792 699984
rect 292540 699944 348792 699972
rect 292540 699932 292546 699944
rect 348786 699932 348792 699944
rect 348844 699932 348850 699984
rect 289722 699864 289728 699916
rect 289780 699904 289786 699916
rect 332502 699904 332508 699916
rect 289780 699876 332508 699904
rect 289780 699864 289786 699876
rect 332502 699864 332508 699876
rect 332560 699864 332566 699916
rect 267642 699796 267648 699848
rect 267700 699836 267706 699848
rect 296714 699836 296720 699848
rect 267700 699808 296720 699836
rect 267700 699796 267706 699808
rect 296714 699796 296720 699808
rect 296772 699796 296778 699848
rect 283834 699728 283840 699780
rect 283892 699768 283898 699780
rect 299566 699768 299572 699780
rect 283892 699740 299572 699768
rect 283892 699728 283898 699740
rect 299566 699728 299572 699740
rect 299624 699728 299630 699780
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 253842 696940 253848 696992
rect 253900 696980 253906 696992
rect 580166 696980 580172 696992
rect 253900 696952 580172 696980
rect 253900 696940 253906 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 256602 683204 256608 683256
rect 256660 683244 256666 683256
rect 580166 683244 580172 683256
rect 256660 683216 580172 683244
rect 256660 683204 256666 683216
rect 580166 683204 580172 683216
rect 580224 683204 580230 683256
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 338114 683176 338120 683188
rect 3476 683148 338120 683176
rect 3476 683136 3482 683148
rect 338114 683136 338120 683148
rect 338172 683136 338178 683188
rect 251082 670760 251088 670812
rect 251140 670800 251146 670812
rect 580166 670800 580172 670812
rect 251140 670772 580172 670800
rect 251140 670760 251146 670772
rect 580166 670760 580172 670772
rect 580224 670760 580230 670812
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 345014 670732 345020 670744
rect 3568 670704 345020 670732
rect 3568 670692 3574 670704
rect 345014 670692 345020 670704
rect 345072 670692 345078 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 340874 656928 340880 656940
rect 3476 656900 340880 656928
rect 3476 656888 3482 656900
rect 340874 656888 340880 656900
rect 340932 656888 340938 656940
rect 244182 643084 244188 643136
rect 244240 643124 244246 643136
rect 580166 643124 580172 643136
rect 244240 643096 580172 643124
rect 244240 643084 244246 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 347774 632108 347780 632120
rect 3476 632080 347780 632108
rect 3476 632068 3482 632080
rect 347774 632068 347780 632080
rect 347832 632068 347838 632120
rect 248322 630640 248328 630692
rect 248380 630680 248386 630692
rect 580166 630680 580172 630692
rect 248380 630652 580172 630680
rect 248380 630640 248386 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 353294 618304 353300 618316
rect 3200 618276 353300 618304
rect 3200 618264 3206 618276
rect 353294 618264 353300 618276
rect 353352 618264 353358 618316
rect 241422 616836 241428 616888
rect 241480 616876 241486 616888
rect 580166 616876 580172 616888
rect 241480 616848 580172 616876
rect 241480 616836 241486 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 350534 605860 350540 605872
rect 3292 605832 350540 605860
rect 3292 605820 3298 605832
rect 350534 605820 350540 605832
rect 350592 605820 350598 605872
rect 235810 590656 235816 590708
rect 235868 590696 235874 590708
rect 579798 590696 579804 590708
rect 235868 590668 579804 590696
rect 235868 590656 235874 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 356054 579680 356060 579692
rect 3384 579652 356060 579680
rect 3384 579640 3390 579652
rect 356054 579640 356060 579652
rect 356112 579640 356118 579692
rect 238662 576852 238668 576904
rect 238720 576892 238726 576904
rect 580166 576892 580172 576904
rect 238720 576864 580172 576892
rect 238720 576852 238726 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 362862 565876 362868 565888
rect 3476 565848 362868 565876
rect 3476 565836 3482 565848
rect 362862 565836 362868 565848
rect 362920 565836 362926 565888
rect 232314 563048 232320 563100
rect 232372 563088 232378 563100
rect 579798 563088 579804 563100
rect 232372 563060 579804 563088
rect 232372 563048 232378 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 247126 561620 247132 561672
rect 247184 561660 247190 561672
rect 248322 561660 248328 561672
rect 247184 561632 248328 561660
rect 247184 561620 247190 561632
rect 248322 561620 248328 561632
rect 248380 561620 248386 561672
rect 250070 561620 250076 561672
rect 250128 561660 250134 561672
rect 251082 561660 251088 561672
rect 250128 561632 251088 561660
rect 250128 561620 250134 561632
rect 251082 561620 251088 561632
rect 251140 561620 251146 561672
rect 253014 561620 253020 561672
rect 253072 561660 253078 561672
rect 253842 561660 253848 561672
rect 253072 561632 253848 561660
rect 253072 561620 253078 561632
rect 253842 561620 253848 561632
rect 253900 561620 253906 561672
rect 270862 561620 270868 561672
rect 270920 561660 270926 561672
rect 271782 561660 271788 561672
rect 270920 561632 271788 561660
rect 270920 561620 270926 561632
rect 271782 561620 271788 561632
rect 271840 561620 271846 561672
rect 273806 561620 273812 561672
rect 273864 561660 273870 561672
rect 274542 561660 274548 561672
rect 273864 561632 274548 561660
rect 273864 561620 273870 561632
rect 274542 561620 274548 561632
rect 274600 561620 274606 561672
rect 288618 561620 288624 561672
rect 288676 561660 288682 561672
rect 289722 561660 289728 561672
rect 288676 561632 289728 561660
rect 288676 561620 288682 561632
rect 289722 561620 289728 561632
rect 289780 561620 289786 561672
rect 291654 561620 291660 561672
rect 291712 561660 291718 561672
rect 292482 561660 292488 561672
rect 291712 561632 292488 561660
rect 291712 561620 291718 561632
rect 292482 561620 292488 561632
rect 292540 561620 292546 561672
rect 294598 561484 294604 561536
rect 294656 561524 294662 561536
rect 299474 561524 299480 561536
rect 294656 561496 299480 561524
rect 294656 561484 294662 561496
rect 299474 561484 299480 561496
rect 299532 561484 299538 561536
rect 235902 561416 235908 561468
rect 235960 561456 235966 561468
rect 303522 561456 303528 561468
rect 235960 561428 303528 561456
rect 235960 561416 235966 561428
rect 303522 561416 303528 561428
rect 303580 561416 303586 561468
rect 285674 561348 285680 561400
rect 285732 561388 285738 561400
rect 364334 561388 364340 561400
rect 285732 561360 364340 561388
rect 285732 561348 285738 561360
rect 364334 561348 364340 561360
rect 364392 561348 364398 561400
rect 171042 561280 171048 561332
rect 171100 561320 171106 561332
rect 312446 561320 312452 561332
rect 171100 561292 312452 561320
rect 171100 561280 171106 561292
rect 312446 561280 312452 561292
rect 312504 561280 312510 561332
rect 276750 561212 276756 561264
rect 276808 561252 276814 561264
rect 429194 561252 429200 561264
rect 276808 561224 429200 561252
rect 276808 561212 276814 561224
rect 429194 561212 429200 561224
rect 429252 561212 429258 561264
rect 106182 561144 106188 561196
rect 106240 561184 106246 561196
rect 321278 561184 321284 561196
rect 106240 561156 321284 561184
rect 106240 561144 106246 561156
rect 321278 561144 321284 561156
rect 321336 561144 321342 561196
rect 267918 561076 267924 561128
rect 267976 561116 267982 561128
rect 494054 561116 494060 561128
rect 267976 561088 494060 561116
rect 267976 561076 267982 561088
rect 494054 561076 494060 561088
rect 494112 561076 494118 561128
rect 211522 561008 211528 561060
rect 211580 561048 211586 561060
rect 486418 561048 486424 561060
rect 211580 561020 486424 561048
rect 211580 561008 211586 561020
rect 486418 561008 486424 561020
rect 486476 561008 486482 561060
rect 258994 560940 259000 560992
rect 259052 560980 259058 560992
rect 558914 560980 558920 560992
rect 259052 560952 558920 560980
rect 259052 560940 259058 560952
rect 558914 560940 558920 560952
rect 558972 560940 558978 560992
rect 202598 560872 202604 560924
rect 202656 560912 202662 560924
rect 485038 560912 485044 560924
rect 202656 560884 485044 560912
rect 202656 560872 202662 560884
rect 485038 560872 485044 560884
rect 485096 560872 485102 560924
rect 193674 560804 193680 560856
rect 193732 560844 193738 560856
rect 483658 560844 483664 560856
rect 193732 560816 483664 560844
rect 193732 560804 193738 560816
rect 483658 560804 483664 560816
rect 483716 560804 483722 560856
rect 184842 560736 184848 560788
rect 184900 560776 184906 560788
rect 482278 560776 482284 560788
rect 184900 560748 482284 560776
rect 184900 560736 184906 560748
rect 482278 560736 482284 560748
rect 482336 560736 482342 560788
rect 175918 560668 175924 560720
rect 175976 560708 175982 560720
rect 479518 560708 479524 560720
rect 175976 560680 479524 560708
rect 175976 560668 175982 560680
rect 479518 560668 479524 560680
rect 479576 560668 479582 560720
rect 166994 560600 167000 560652
rect 167052 560640 167058 560652
rect 475378 560640 475384 560652
rect 167052 560612 475384 560640
rect 167052 560600 167058 560612
rect 475378 560600 475384 560612
rect 475436 560600 475442 560652
rect 29638 560532 29644 560584
rect 29696 560572 29702 560584
rect 398466 560572 398472 560584
rect 29696 560544 398472 560572
rect 29696 560532 29702 560544
rect 398466 560532 398472 560544
rect 398524 560532 398530 560584
rect 32398 560464 32404 560516
rect 32456 560504 32462 560516
rect 407390 560504 407396 560516
rect 32456 560476 407396 560504
rect 32456 560464 32462 560476
rect 407390 560464 407396 560476
rect 407448 560464 407454 560516
rect 33778 560396 33784 560448
rect 33836 560436 33842 560448
rect 416222 560436 416228 560448
rect 33836 560408 416228 560436
rect 33836 560396 33842 560408
rect 416222 560396 416228 560408
rect 416280 560396 416286 560448
rect 35158 560328 35164 560380
rect 35216 560368 35222 560380
rect 425146 560368 425152 560380
rect 35216 560340 425152 560368
rect 35216 560328 35222 560340
rect 425146 560328 425152 560340
rect 425204 560328 425210 560380
rect 36538 560260 36544 560312
rect 36596 560300 36602 560312
rect 434070 560300 434076 560312
rect 36596 560272 434076 560300
rect 36596 560260 36602 560272
rect 434070 560260 434076 560272
rect 434128 560260 434134 560312
rect 205542 559580 205548 559632
rect 205600 559620 205606 559632
rect 468478 559620 468484 559632
rect 205600 559592 468484 559620
rect 205600 559580 205606 559592
rect 468478 559580 468484 559592
rect 468536 559580 468542 559632
rect 115198 559512 115204 559564
rect 115256 559552 115262 559564
rect 380618 559552 380624 559564
rect 115256 559524 380624 559552
rect 115256 559512 115262 559524
rect 380618 559512 380624 559524
rect 380676 559512 380682 559564
rect 196710 559444 196716 559496
rect 196768 559484 196774 559496
rect 467098 559484 467104 559496
rect 196768 559456 467104 559484
rect 196768 559444 196774 559456
rect 467098 559444 467104 559456
rect 467156 559444 467162 559496
rect 122098 559376 122104 559428
rect 122156 559416 122162 559428
rect 395522 559416 395528 559428
rect 122156 559388 395528 559416
rect 122156 559376 122162 559388
rect 395522 559376 395528 559388
rect 395580 559376 395586 559428
rect 190730 559308 190736 559360
rect 190788 559348 190794 559360
rect 497458 559348 497464 559360
rect 190788 559320 497464 559348
rect 190788 559308 190794 559320
rect 497458 559308 497464 559320
rect 497516 559308 497522 559360
rect 108298 559240 108304 559292
rect 108356 559280 108362 559292
rect 422202 559280 422208 559292
rect 108356 559252 422208 559280
rect 108356 559240 108362 559252
rect 422202 559240 422208 559252
rect 422260 559240 422266 559292
rect 172974 559172 172980 559224
rect 173032 559212 173038 559224
rect 490558 559212 490564 559224
rect 173032 559184 490564 559212
rect 173032 559172 173038 559184
rect 490558 559172 490564 559184
rect 490616 559172 490622 559224
rect 155126 559104 155132 559156
rect 155184 559144 155190 559156
rect 472618 559144 472624 559156
rect 155184 559116 472624 559144
rect 155184 559104 155190 559116
rect 472618 559104 472624 559116
rect 472676 559104 472682 559156
rect 83458 559036 83464 559088
rect 83516 559076 83522 559088
rect 428090 559076 428096 559088
rect 83516 559048 428096 559076
rect 83516 559036 83522 559048
rect 428090 559036 428096 559048
rect 428148 559036 428154 559088
rect 169938 558968 169944 559020
rect 169996 559008 170002 559020
rect 522298 559008 522304 559020
rect 169996 558980 522304 559008
rect 169996 558968 170002 558980
rect 522298 558968 522304 558980
rect 522356 558968 522362 559020
rect 4798 558900 4804 558952
rect 4856 558940 4862 558952
rect 410334 558940 410340 558952
rect 4856 558912 410340 558940
rect 4856 558900 4862 558912
rect 410334 558900 410340 558912
rect 410392 558900 410398 558952
rect 214466 558220 214472 558272
rect 214524 558260 214530 558272
rect 462958 558260 462964 558272
rect 214524 558232 462964 558260
rect 214524 558220 214530 558232
rect 462958 558220 462964 558232
rect 463016 558220 463022 558272
rect 187786 558152 187792 558204
rect 187844 558192 187850 558204
rect 465718 558192 465724 558204
rect 187844 558164 465724 558192
rect 187844 558152 187850 558164
rect 465718 558152 465724 558164
rect 465776 558152 465782 558204
rect 178862 558084 178868 558136
rect 178920 558124 178926 558136
rect 464338 558124 464344 558136
rect 178920 558096 464344 558124
rect 178920 558084 178926 558096
rect 464338 558084 464344 558096
rect 464396 558084 464402 558136
rect 123478 558016 123484 558068
rect 123536 558056 123542 558068
rect 412910 558056 412916 558068
rect 123536 558028 412916 558056
rect 123536 558016 123542 558028
rect 412910 558016 412916 558028
rect 412968 558016 412974 558068
rect 199838 557948 199844 558000
rect 199896 557988 199902 558000
rect 500218 557988 500224 558000
rect 199896 557960 500224 557988
rect 199896 557948 199902 557960
rect 500218 557948 500224 557960
rect 500276 557948 500282 558000
rect 79318 557880 79324 557932
rect 79376 557920 79382 557932
rect 386414 557920 386420 557932
rect 79376 557892 386420 557920
rect 79376 557880 79382 557892
rect 386414 557880 386420 557892
rect 386472 557880 386478 557932
rect 119338 557812 119344 557864
rect 119396 557852 119402 557864
rect 430758 557852 430764 557864
rect 119396 557824 430764 557852
rect 119396 557812 119402 557824
rect 430758 557812 430764 557824
rect 430816 557812 430822 557864
rect 182082 557744 182088 557796
rect 182140 557784 182146 557796
rect 493318 557784 493324 557796
rect 182140 557756 493324 557784
rect 182140 557744 182146 557756
rect 493318 557744 493324 557756
rect 493376 557744 493382 557796
rect 164142 557676 164148 557728
rect 164200 557716 164206 557728
rect 489178 557716 489184 557728
rect 164200 557688 489184 557716
rect 164200 557676 164206 557688
rect 489178 557676 489184 557688
rect 489236 557676 489242 557728
rect 128722 557608 128728 557660
rect 128780 557648 128786 557660
rect 471238 557648 471244 557660
rect 128780 557620 471244 557648
rect 128780 557608 128786 557620
rect 471238 557608 471244 557620
rect 471296 557608 471302 557660
rect 11698 557540 11704 557592
rect 11756 557580 11762 557592
rect 418982 557580 418988 557592
rect 11756 557552 418988 557580
rect 11756 557540 11762 557552
rect 418982 557540 418988 557552
rect 419040 557540 419046 557592
rect 359550 557444 359556 557456
rect 219406 557416 223620 557444
rect 359511 557416 359556 557444
rect 161290 557376 161296 557388
rect 161251 557348 161296 557376
rect 161290 557336 161296 557348
rect 161348 557336 161354 557388
rect 208946 557376 208952 557388
rect 208907 557348 208952 557376
rect 208946 557336 208952 557348
rect 209004 557336 209010 557388
rect 217778 557376 217784 557388
rect 217739 557348 217784 557376
rect 217778 557336 217784 557348
rect 217836 557336 217842 557388
rect 3326 557200 3332 557252
rect 3384 557240 3390 557252
rect 219406 557240 219434 557416
rect 220722 557336 220728 557388
rect 220780 557336 220786 557388
rect 223482 557336 223488 557388
rect 223540 557336 223546 557388
rect 3384 557212 219434 557240
rect 3384 557200 3390 557212
rect 220740 557104 220768 557336
rect 223500 557172 223528 557336
rect 223592 557240 223620 557416
rect 359550 557404 359556 557416
rect 359608 557404 359614 557456
rect 365622 557444 365628 557456
rect 365583 557416 365628 557444
rect 365622 557404 365628 557416
rect 365680 557404 365686 557456
rect 368474 557444 368480 557456
rect 368435 557416 368480 557444
rect 368474 557404 368480 557416
rect 368532 557404 368538 557456
rect 371510 557444 371516 557456
rect 371471 557416 371516 557444
rect 371510 557404 371516 557416
rect 371568 557404 371574 557456
rect 374454 557444 374460 557456
rect 374415 557416 374460 557444
rect 374454 557404 374460 557416
rect 374512 557404 374518 557456
rect 377398 557444 377404 557456
rect 377359 557416 377404 557444
rect 377398 557404 377404 557416
rect 377456 557404 377462 557456
rect 383746 557444 383752 557456
rect 383707 557416 383752 557444
rect 383746 557404 383752 557416
rect 383804 557404 383810 557456
rect 389174 557444 389180 557456
rect 389135 557416 389180 557444
rect 389174 557404 389180 557416
rect 389232 557404 389238 557456
rect 392118 557444 392124 557456
rect 392079 557416 392124 557444
rect 392118 557404 392124 557416
rect 392176 557404 392182 557456
rect 401134 557444 401140 557456
rect 401095 557416 401140 557444
rect 401134 557404 401140 557416
rect 401192 557404 401198 557456
rect 404170 557444 404176 557456
rect 404131 557416 404176 557444
rect 404170 557404 404176 557416
rect 404228 557404 404234 557456
rect 226610 557336 226616 557388
rect 226668 557376 226674 557388
rect 226668 557348 229094 557376
rect 226668 557336 226674 557348
rect 229066 557308 229094 557348
rect 229554 557336 229560 557388
rect 229612 557376 229618 557388
rect 580718 557376 580724 557388
rect 229612 557348 580724 557376
rect 229612 557336 229618 557348
rect 580718 557336 580724 557348
rect 580776 557336 580782 557388
rect 580810 557308 580816 557320
rect 229066 557280 580816 557308
rect 580810 557268 580816 557280
rect 580868 557268 580874 557320
rect 359553 557243 359611 557249
rect 359553 557240 359565 557243
rect 223592 557212 359565 557240
rect 359553 557209 359565 557212
rect 359599 557209 359611 557243
rect 359553 557203 359611 557209
rect 580626 557172 580632 557184
rect 223500 557144 580632 557172
rect 580626 557132 580632 557144
rect 580684 557132 580690 557184
rect 580442 557104 580448 557116
rect 220740 557076 580448 557104
rect 580442 557064 580448 557076
rect 580500 557064 580506 557116
rect 3142 556996 3148 557048
rect 3200 557036 3206 557048
rect 365625 557039 365683 557045
rect 365625 557036 365637 557039
rect 3200 557008 365637 557036
rect 3200 556996 3206 557008
rect 365625 557005 365637 557008
rect 365671 557005 365683 557039
rect 365625 556999 365683 557005
rect 217781 556971 217839 556977
rect 217781 556937 217793 556971
rect 217827 556968 217839 556971
rect 580534 556968 580540 556980
rect 217827 556940 580540 556968
rect 217827 556937 217839 556940
rect 217781 556931 217839 556937
rect 580534 556928 580540 556940
rect 580592 556928 580598 556980
rect 4062 556860 4068 556912
rect 4120 556900 4126 556912
rect 368477 556903 368535 556909
rect 368477 556900 368489 556903
rect 4120 556872 368489 556900
rect 4120 556860 4126 556872
rect 368477 556869 368489 556872
rect 368523 556869 368535 556903
rect 368477 556863 368535 556869
rect 3234 556792 3240 556844
rect 3292 556832 3298 556844
rect 371513 556835 371571 556841
rect 371513 556832 371525 556835
rect 3292 556804 371525 556832
rect 3292 556792 3298 556804
rect 371513 556801 371525 556804
rect 371559 556801 371571 556835
rect 371513 556795 371571 556801
rect 3970 556724 3976 556776
rect 4028 556764 4034 556776
rect 374457 556767 374515 556773
rect 374457 556764 374469 556767
rect 4028 556736 374469 556764
rect 4028 556724 4034 556736
rect 374457 556733 374469 556736
rect 374503 556733 374515 556767
rect 374457 556727 374515 556733
rect 208949 556699 209007 556705
rect 208949 556665 208961 556699
rect 208995 556696 209007 556699
rect 580350 556696 580356 556708
rect 208995 556668 580356 556696
rect 208995 556665 209007 556668
rect 208949 556659 209007 556665
rect 580350 556656 580356 556668
rect 580408 556656 580414 556708
rect 3878 556588 3884 556640
rect 3936 556628 3942 556640
rect 377401 556631 377459 556637
rect 377401 556628 377413 556631
rect 3936 556600 377413 556628
rect 3936 556588 3942 556600
rect 377401 556597 377413 556600
rect 377447 556597 377459 556631
rect 377401 556591 377459 556597
rect 3786 556520 3792 556572
rect 3844 556560 3850 556572
rect 383749 556563 383807 556569
rect 383749 556560 383761 556563
rect 3844 556532 383761 556560
rect 3844 556520 3850 556532
rect 383749 556529 383761 556532
rect 383795 556529 383807 556563
rect 383749 556523 383807 556529
rect 3694 556452 3700 556504
rect 3752 556492 3758 556504
rect 389177 556495 389235 556501
rect 389177 556492 389189 556495
rect 3752 556464 389189 556492
rect 3752 556452 3758 556464
rect 389177 556461 389189 556464
rect 389223 556461 389235 556495
rect 389177 556455 389235 556461
rect 3602 556384 3608 556436
rect 3660 556424 3666 556436
rect 392121 556427 392179 556433
rect 392121 556424 392133 556427
rect 3660 556396 392133 556424
rect 3660 556384 3666 556396
rect 392121 556393 392133 556396
rect 392167 556393 392179 556427
rect 392121 556387 392179 556393
rect 3510 556316 3516 556368
rect 3568 556356 3574 556368
rect 401137 556359 401195 556365
rect 401137 556356 401149 556359
rect 3568 556328 401149 556356
rect 3568 556316 3574 556328
rect 401137 556325 401149 556328
rect 401183 556325 401195 556359
rect 401137 556319 401195 556325
rect 3418 556248 3424 556300
rect 3476 556288 3482 556300
rect 404173 556291 404231 556297
rect 404173 556288 404185 556291
rect 3476 556260 404185 556288
rect 3476 556248 3482 556260
rect 404173 556257 404185 556260
rect 404219 556257 404231 556291
rect 404173 556251 404231 556257
rect 161293 556223 161351 556229
rect 161293 556189 161305 556223
rect 161339 556220 161351 556223
rect 580258 556220 580264 556232
rect 161339 556192 580264 556220
rect 161339 556189 161351 556192
rect 161293 556183 161351 556189
rect 580258 556180 580264 556192
rect 580316 556180 580322 556232
rect 2866 463632 2872 463684
rect 2924 463672 2930 463684
rect 115198 463672 115204 463684
rect 2924 463644 115204 463672
rect 2924 463632 2930 463644
rect 115198 463632 115204 463644
rect 115256 463632 115262 463684
rect 462958 458124 462964 458176
rect 463016 458164 463022 458176
rect 580166 458164 580172 458176
rect 463016 458136 580172 458164
rect 463016 458124 463022 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 486418 419432 486424 419484
rect 486476 419472 486482 419484
rect 580166 419472 580172 419484
rect 486476 419444 580172 419472
rect 486476 419432 486482 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 468478 405628 468484 405680
rect 468536 405668 468542 405680
rect 579614 405668 579620 405680
rect 468536 405640 579620 405668
rect 468536 405628 468542 405640
rect 579614 405628 579620 405640
rect 579672 405628 579678 405680
rect 3326 398760 3332 398812
rect 3384 398800 3390 398812
rect 79318 398800 79324 398812
rect 3384 398772 79324 398800
rect 3384 398760 3390 398772
rect 79318 398760 79324 398772
rect 79376 398760 79382 398812
rect 500218 379448 500224 379500
rect 500276 379488 500282 379500
rect 580166 379488 580172 379500
rect 500276 379460 580172 379488
rect 500276 379448 500282 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 485038 365644 485044 365696
rect 485096 365684 485102 365696
rect 580166 365684 580172 365696
rect 485096 365656 580172 365684
rect 485096 365644 485102 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 29638 358748 29644 358760
rect 3384 358720 29644 358748
rect 3384 358708 3390 358720
rect 29638 358708 29644 358720
rect 29696 358708 29702 358760
rect 467098 353200 467104 353252
rect 467156 353240 467162 353252
rect 580166 353240 580172 353252
rect 467156 353212 580172 353240
rect 467156 353200 467162 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3326 346332 3332 346384
rect 3384 346372 3390 346384
rect 122098 346372 122104 346384
rect 3384 346344 122104 346372
rect 3384 346332 3390 346344
rect 122098 346332 122104 346344
rect 122156 346332 122162 346384
rect 497458 325592 497464 325644
rect 497516 325632 497522 325644
rect 579890 325632 579896 325644
rect 497516 325604 579896 325632
rect 497516 325592 497522 325604
rect 579890 325592 579896 325604
rect 579948 325592 579954 325644
rect 483658 313216 483664 313268
rect 483716 313256 483722 313268
rect 580166 313256 580172 313268
rect 483716 313228 580172 313256
rect 483716 313216 483722 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3510 306280 3516 306332
rect 3568 306320 3574 306332
rect 32398 306320 32404 306332
rect 3568 306292 32404 306320
rect 3568 306280 3574 306292
rect 32398 306280 32404 306292
rect 32456 306280 32462 306332
rect 465718 299412 465724 299464
rect 465776 299452 465782 299464
rect 579614 299452 579620 299464
rect 465776 299424 579620 299452
rect 465776 299412 465782 299424
rect 579614 299412 579620 299424
rect 579672 299412 579678 299464
rect 493318 273164 493324 273216
rect 493376 273204 493382 273216
rect 579890 273204 579896 273216
rect 493376 273176 579896 273204
rect 493376 273164 493382 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 2774 267384 2780 267436
rect 2832 267424 2838 267436
rect 4798 267424 4804 267436
rect 2832 267396 4804 267424
rect 2832 267384 2838 267396
rect 4798 267384 4804 267396
rect 4856 267384 4862 267436
rect 482278 259360 482284 259412
rect 482336 259400 482342 259412
rect 579798 259400 579804 259412
rect 482336 259372 579804 259400
rect 482336 259360 482342 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 3418 255212 3424 255264
rect 3476 255252 3482 255264
rect 33778 255252 33784 255264
rect 3476 255224 33784 255252
rect 3476 255212 3482 255224
rect 33778 255212 33784 255224
rect 33836 255212 33842 255264
rect 464338 245556 464344 245608
rect 464396 245596 464402 245608
rect 580166 245596 580172 245608
rect 464396 245568 580172 245596
rect 464396 245556 464402 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3418 241408 3424 241460
rect 3476 241448 3482 241460
rect 123478 241448 123484 241460
rect 3476 241420 123484 241448
rect 3476 241408 3482 241420
rect 123478 241408 123484 241420
rect 123536 241408 123542 241460
rect 490558 233180 490564 233232
rect 490616 233220 490622 233232
rect 580166 233220 580172 233232
rect 490616 233192 580172 233220
rect 490616 233180 490622 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 479518 219376 479524 219428
rect 479576 219416 479582 219428
rect 579890 219416 579896 219428
rect 479576 219388 579896 219416
rect 479576 219376 479582 219388
rect 579890 219376 579896 219388
rect 579948 219376 579954 219428
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 11698 215268 11704 215280
rect 3384 215240 11704 215268
rect 3384 215228 3390 215240
rect 11698 215228 11704 215240
rect 11756 215228 11762 215280
rect 522298 206932 522304 206984
rect 522356 206972 522362 206984
rect 580166 206972 580172 206984
rect 522356 206944 580172 206972
rect 522356 206932 522362 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 3418 202784 3424 202836
rect 3476 202824 3482 202836
rect 35158 202824 35164 202836
rect 3476 202796 35164 202824
rect 3476 202784 3482 202796
rect 35158 202784 35164 202796
rect 35216 202784 35222 202836
rect 489178 193128 489184 193180
rect 489236 193168 489242 193180
rect 580166 193168 580172 193180
rect 489236 193140 580172 193168
rect 489236 193128 489242 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 108298 189020 108304 189032
rect 3476 188992 108304 189020
rect 3476 188980 3482 188992
rect 108298 188980 108304 188992
rect 108356 188980 108362 189032
rect 475378 179324 475384 179376
rect 475436 179364 475442 179376
rect 579982 179364 579988 179376
rect 475436 179336 579988 179364
rect 475436 179324 475442 179336
rect 579982 179324 579988 179336
rect 580040 179324 580046 179376
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 83458 164200 83464 164212
rect 3292 164172 83464 164200
rect 3292 164160 3298 164172
rect 83458 164160 83464 164172
rect 83516 164160 83522 164212
rect 472618 153144 472624 153196
rect 472676 153184 472682 153196
rect 580166 153184 580172 153196
rect 472676 153156 580172 153184
rect 472676 153144 472682 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 36538 150396 36544 150408
rect 3476 150368 36544 150396
rect 3476 150356 3482 150368
rect 36538 150356 36544 150368
rect 36596 150356 36602 150408
rect 107562 148996 107568 149048
rect 107620 149036 107626 149048
rect 186038 149036 186044 149048
rect 107620 149008 186044 149036
rect 107620 148996 107626 149008
rect 186038 148996 186044 149008
rect 186096 148996 186102 149048
rect 191742 148996 191748 149048
rect 191800 149036 191806 149048
rect 234706 149036 234712 149048
rect 191800 149008 234712 149036
rect 191800 148996 191806 149008
rect 234706 148996 234712 149008
rect 234764 148996 234770 149048
rect 241422 148996 241428 149048
rect 241480 149036 241486 149048
rect 263594 149036 263600 149048
rect 241480 149008 263600 149036
rect 241480 148996 241486 149008
rect 263594 148996 263600 149008
rect 263652 148996 263658 149048
rect 270402 148996 270408 149048
rect 270460 149036 270466 149048
rect 280706 149036 280712 149048
rect 270460 149008 280712 149036
rect 270460 148996 270466 149008
rect 280706 148996 280712 149008
rect 280764 148996 280770 149048
rect 372614 148996 372620 149048
rect 372672 149036 372678 149048
rect 374638 149036 374644 149048
rect 372672 149008 374644 149036
rect 372672 148996 372678 149008
rect 374638 148996 374644 149008
rect 374696 148996 374702 149048
rect 406286 148996 406292 149048
rect 406344 149036 406350 149048
rect 485774 149036 485780 149048
rect 406344 149008 485780 149036
rect 406344 148996 406350 149008
rect 485774 148996 485780 149008
rect 485832 148996 485838 149048
rect 104158 148928 104164 148980
rect 104216 148968 104222 148980
rect 183278 148968 183284 148980
rect 104216 148940 183284 148968
rect 104216 148928 104222 148940
rect 183278 148928 183284 148940
rect 183336 148928 183342 148980
rect 187602 148928 187608 148980
rect 187660 148968 187666 148980
rect 232682 148968 232688 148980
rect 187660 148940 232688 148968
rect 187660 148928 187666 148940
rect 232682 148928 232688 148940
rect 232740 148928 232746 148980
rect 235902 148928 235908 148980
rect 235960 148968 235966 148980
rect 260098 148968 260104 148980
rect 235960 148940 260104 148968
rect 235960 148928 235966 148940
rect 260098 148928 260104 148940
rect 260156 148928 260162 148980
rect 260742 148928 260748 148980
rect 260800 148968 260806 148980
rect 274542 148968 274548 148980
rect 260800 148940 274548 148968
rect 260800 148928 260806 148940
rect 274542 148928 274548 148940
rect 274600 148928 274606 148980
rect 347958 148928 347964 148980
rect 348016 148968 348022 148980
rect 385218 148968 385224 148980
rect 348016 148940 385224 148968
rect 348016 148928 348022 148940
rect 385218 148928 385224 148940
rect 385276 148928 385282 148980
rect 410426 148928 410432 148980
rect 410484 148968 410490 148980
rect 492674 148968 492680 148980
rect 410484 148940 492680 148968
rect 410484 148928 410490 148940
rect 492674 148928 492680 148940
rect 492732 148928 492738 148980
rect 93118 148860 93124 148912
rect 93176 148900 93182 148912
rect 177114 148900 177120 148912
rect 93176 148872 177120 148900
rect 93176 148860 93182 148872
rect 177114 148860 177120 148872
rect 177172 148860 177178 148912
rect 177298 148860 177304 148912
rect 177356 148900 177362 148912
rect 181254 148900 181260 148912
rect 177356 148872 181260 148900
rect 177356 148860 177362 148872
rect 181254 148860 181260 148872
rect 181312 148860 181318 148912
rect 184198 148860 184204 148912
rect 184256 148900 184262 148912
rect 229922 148900 229928 148912
rect 184256 148872 229928 148900
rect 184256 148860 184262 148872
rect 229922 148860 229928 148872
rect 229980 148860 229986 148912
rect 238662 148860 238668 148912
rect 238720 148900 238726 148912
rect 262214 148900 262220 148912
rect 238720 148872 262220 148900
rect 238720 148860 238726 148872
rect 262214 148860 262220 148872
rect 262272 148860 262278 148912
rect 264882 148860 264888 148912
rect 264940 148900 264946 148912
rect 276934 148900 276940 148912
rect 264940 148872 276940 148900
rect 264940 148860 264946 148872
rect 276934 148860 276940 148872
rect 276992 148860 276998 148912
rect 277210 148860 277216 148912
rect 277268 148900 277274 148912
rect 284110 148900 284116 148912
rect 277268 148872 284116 148900
rect 277268 148860 277274 148872
rect 284110 148860 284116 148872
rect 284168 148860 284174 148912
rect 349338 148860 349344 148912
rect 349396 148900 349402 148912
rect 388070 148900 388076 148912
rect 349396 148872 388076 148900
rect 349396 148860 349402 148872
rect 388070 148860 388076 148872
rect 388128 148860 388134 148912
rect 419994 148860 420000 148912
rect 420052 148900 420058 148912
rect 504358 148900 504364 148912
rect 420052 148872 504364 148900
rect 420052 148860 420058 148872
rect 504358 148860 504364 148872
rect 504416 148860 504422 148912
rect 75178 148792 75184 148844
rect 75236 148832 75242 148844
rect 166810 148832 166816 148844
rect 75236 148804 166816 148832
rect 75236 148792 75242 148804
rect 166810 148792 166816 148804
rect 166868 148792 166874 148844
rect 173158 148792 173164 148844
rect 173216 148832 173222 148844
rect 223758 148832 223764 148844
rect 173216 148804 223764 148832
rect 173216 148792 173222 148804
rect 223758 148792 223764 148804
rect 223816 148792 223822 148844
rect 237282 148792 237288 148844
rect 237340 148832 237346 148844
rect 261478 148832 261484 148844
rect 237340 148804 261484 148832
rect 237340 148792 237346 148804
rect 261478 148792 261484 148804
rect 261536 148792 261542 148844
rect 262858 148792 262864 148844
rect 262916 148832 262922 148844
rect 275922 148832 275928 148844
rect 262916 148804 275928 148832
rect 262916 148792 262922 148804
rect 275922 148792 275928 148804
rect 275980 148792 275986 148844
rect 351362 148792 351368 148844
rect 351420 148832 351426 148844
rect 389726 148832 389732 148844
rect 351420 148804 389732 148832
rect 351420 148792 351426 148804
rect 389726 148792 389732 148804
rect 389784 148792 389790 148844
rect 413094 148792 413100 148844
rect 413152 148832 413158 148844
rect 497458 148832 497464 148844
rect 413152 148804 497464 148832
rect 413152 148792 413158 148804
rect 497458 148792 497464 148804
rect 497516 148792 497522 148844
rect 35158 148724 35164 148776
rect 35216 148764 35222 148776
rect 135254 148764 135260 148776
rect 35216 148736 135260 148764
rect 35216 148724 35222 148736
rect 135254 148724 135260 148736
rect 135312 148724 135318 148776
rect 154850 148724 154856 148776
rect 154908 148764 154914 148776
rect 157886 148764 157892 148776
rect 154908 148736 157892 148764
rect 154908 148724 154914 148736
rect 157886 148724 157892 148736
rect 157944 148724 157950 148776
rect 166258 148724 166264 148776
rect 166316 148764 166322 148776
rect 218974 148764 218980 148776
rect 166316 148736 218980 148764
rect 166316 148724 166322 148736
rect 218974 148724 218980 148736
rect 219032 148724 219038 148776
rect 234522 148724 234528 148776
rect 234580 148764 234586 148776
rect 259454 148764 259460 148776
rect 234580 148736 259460 148764
rect 234580 148724 234586 148736
rect 259454 148724 259460 148736
rect 259512 148724 259518 148776
rect 263502 148724 263508 148776
rect 263560 148764 263566 148776
rect 276566 148764 276572 148776
rect 263560 148736 276572 148764
rect 263560 148724 263566 148736
rect 276566 148724 276572 148736
rect 276624 148724 276630 148776
rect 276658 148724 276664 148776
rect 276716 148764 276722 148776
rect 283466 148764 283472 148776
rect 276716 148736 283472 148764
rect 276716 148724 276722 148736
rect 283466 148724 283472 148736
rect 283524 148724 283530 148776
rect 352742 148724 352748 148776
rect 352800 148764 352806 148776
rect 393498 148764 393504 148776
rect 352800 148736 393504 148764
rect 352800 148724 352806 148736
rect 393498 148724 393504 148736
rect 393556 148724 393562 148776
rect 414474 148724 414480 148776
rect 414532 148764 414538 148776
rect 499574 148764 499580 148776
rect 414532 148736 499580 148764
rect 414532 148724 414538 148736
rect 499574 148724 499580 148736
rect 499632 148724 499638 148776
rect 22738 148656 22744 148708
rect 22796 148696 22802 148708
rect 124950 148696 124956 148708
rect 22796 148668 124956 148696
rect 22796 148656 22802 148668
rect 124950 148656 124956 148668
rect 125008 148656 125014 148708
rect 155218 148656 155224 148708
rect 155276 148696 155282 148708
rect 213454 148696 213460 148708
rect 155276 148668 213460 148696
rect 155276 148656 155282 148668
rect 213454 148656 213460 148668
rect 213512 148656 213518 148708
rect 231762 148656 231768 148708
rect 231820 148696 231826 148708
rect 258074 148696 258080 148708
rect 231820 148668 258080 148696
rect 231820 148656 231826 148668
rect 258074 148656 258080 148668
rect 258132 148656 258138 148708
rect 259362 148656 259368 148708
rect 259420 148696 259426 148708
rect 273806 148696 273812 148708
rect 259420 148668 273812 148696
rect 259420 148656 259426 148668
rect 273806 148656 273812 148668
rect 273864 148656 273870 148708
rect 274542 148656 274548 148708
rect 274600 148696 274606 148708
rect 282730 148696 282736 148708
rect 274600 148668 282736 148696
rect 274600 148656 274606 148668
rect 282730 148656 282736 148668
rect 282788 148656 282794 148708
rect 356882 148656 356888 148708
rect 356940 148696 356946 148708
rect 400398 148696 400404 148708
rect 356940 148668 400404 148696
rect 356940 148656 356946 148668
rect 400398 148656 400404 148668
rect 400456 148656 400462 148708
rect 409046 148656 409052 148708
rect 409104 148696 409110 148708
rect 410794 148696 410800 148708
rect 409104 148668 410800 148696
rect 409104 148656 409110 148668
rect 410794 148656 410800 148668
rect 410852 148656 410858 148708
rect 417234 148656 417240 148708
rect 417292 148696 417298 148708
rect 502978 148696 502984 148708
rect 417292 148668 502984 148696
rect 417292 148656 417298 148668
rect 502978 148656 502984 148668
rect 503036 148656 503042 148708
rect 25498 148588 25504 148640
rect 25556 148628 25562 148640
rect 131850 148628 131856 148640
rect 25556 148600 131856 148628
rect 25556 148588 25562 148600
rect 131850 148588 131856 148600
rect 131908 148588 131914 148640
rect 144362 148588 144368 148640
rect 144420 148628 144426 148640
rect 203150 148628 203156 148640
rect 144420 148600 203156 148628
rect 144420 148588 144426 148600
rect 203150 148588 203156 148600
rect 203208 148588 203214 148640
rect 227622 148588 227628 148640
rect 227680 148628 227686 148640
rect 256050 148628 256056 148640
rect 227680 148600 256056 148628
rect 227680 148588 227686 148600
rect 256050 148588 256056 148600
rect 256108 148588 256114 148640
rect 260650 148588 260656 148640
rect 260708 148628 260714 148640
rect 275186 148628 275192 148640
rect 260708 148600 275192 148628
rect 260708 148588 260714 148600
rect 275186 148588 275192 148600
rect 275244 148588 275250 148640
rect 277302 148588 277308 148640
rect 277360 148628 277366 148640
rect 284846 148628 284852 148640
rect 277360 148600 284852 148628
rect 277360 148588 277366 148600
rect 284846 148588 284852 148600
rect 284904 148588 284910 148640
rect 370590 148588 370596 148640
rect 370648 148628 370654 148640
rect 414658 148628 414664 148640
rect 370648 148600 414664 148628
rect 370648 148588 370654 148600
rect 414658 148588 414664 148600
rect 414716 148588 414722 148640
rect 418614 148588 418620 148640
rect 418672 148628 418678 148640
rect 506474 148628 506480 148640
rect 418672 148600 506480 148628
rect 418672 148588 418678 148600
rect 506474 148588 506480 148600
rect 506532 148588 506538 148640
rect 14458 148520 14464 148572
rect 14516 148560 14522 148572
rect 124306 148560 124312 148572
rect 14516 148532 124312 148560
rect 14516 148520 14522 148532
rect 124306 148520 124312 148532
rect 124364 148520 124370 148572
rect 147122 148520 147128 148572
rect 147180 148560 147186 148572
rect 207290 148560 207296 148572
rect 147180 148532 207296 148560
rect 147180 148520 147186 148532
rect 207290 148520 207296 148532
rect 207348 148520 207354 148572
rect 223482 148520 223488 148572
rect 223540 148560 223546 148572
rect 253290 148560 253296 148572
rect 223540 148532 253296 148560
rect 223540 148520 223546 148532
rect 253290 148520 253296 148532
rect 253348 148520 253354 148572
rect 253842 148520 253848 148572
rect 253900 148560 253906 148572
rect 271138 148560 271144 148572
rect 253900 148532 271144 148560
rect 253900 148520 253906 148532
rect 271138 148520 271144 148532
rect 271196 148520 271202 148572
rect 271782 148520 271788 148572
rect 271840 148560 271846 148572
rect 281350 148560 281356 148572
rect 271840 148532 281356 148560
rect 271840 148520 271846 148532
rect 281350 148520 281356 148532
rect 281408 148520 281414 148572
rect 328730 148520 328736 148572
rect 328788 148560 328794 148572
rect 352006 148560 352012 148572
rect 328788 148532 352012 148560
rect 328788 148520 328794 148532
rect 352006 148520 352012 148532
rect 352064 148520 352070 148572
rect 356146 148520 356152 148572
rect 356204 148560 356210 148572
rect 357342 148560 357348 148572
rect 356204 148532 357348 148560
rect 356204 148520 356210 148532
rect 357342 148520 357348 148532
rect 357400 148520 357406 148572
rect 360286 148520 360292 148572
rect 360344 148560 360350 148572
rect 406378 148560 406384 148572
rect 360344 148532 406384 148560
rect 360344 148520 360350 148532
rect 406378 148520 406384 148532
rect 406436 148520 406442 148572
rect 422754 148520 422760 148572
rect 422812 148560 422818 148572
rect 514754 148560 514760 148572
rect 422812 148532 514760 148560
rect 422812 148520 422818 148532
rect 514754 148520 514760 148532
rect 514812 148520 514818 148572
rect 18598 148452 18604 148504
rect 18656 148492 18662 148504
rect 133138 148492 133144 148504
rect 18656 148464 133144 148492
rect 18656 148452 18662 148464
rect 133138 148452 133144 148464
rect 133196 148452 133202 148504
rect 133322 148452 133328 148504
rect 133380 148492 133386 148504
rect 199010 148492 199016 148504
rect 133380 148464 199016 148492
rect 133380 148452 133386 148464
rect 199010 148452 199016 148464
rect 199068 148452 199074 148504
rect 224862 148452 224868 148504
rect 224920 148492 224926 148504
rect 253934 148492 253940 148504
rect 224920 148464 253940 148492
rect 224920 148452 224926 148464
rect 253934 148452 253940 148464
rect 253992 148452 253998 148504
rect 256602 148452 256608 148504
rect 256660 148492 256666 148504
rect 272518 148492 272524 148504
rect 256660 148464 272524 148492
rect 256660 148452 256666 148464
rect 272518 148452 272524 148464
rect 272576 148452 272582 148504
rect 273898 148452 273904 148504
rect 273956 148492 273962 148504
rect 282086 148492 282092 148504
rect 273956 148464 282092 148492
rect 273956 148452 273962 148464
rect 282086 148452 282092 148464
rect 282144 148452 282150 148504
rect 322566 148452 322572 148504
rect 322624 148492 322630 148504
rect 338758 148492 338764 148504
rect 322624 148464 338764 148492
rect 322624 148452 322630 148464
rect 338758 148452 338764 148464
rect 338816 148452 338822 148504
rect 347222 148452 347228 148504
rect 347280 148492 347286 148504
rect 377398 148492 377404 148504
rect 347280 148464 377404 148492
rect 347280 148452 347286 148464
rect 377398 148452 377404 148464
rect 377456 148452 377462 148504
rect 378870 148452 378876 148504
rect 378928 148492 378934 148504
rect 425698 148492 425704 148504
rect 378928 148464 425704 148492
rect 378928 148452 378934 148464
rect 425698 148452 425704 148464
rect 425756 148452 425762 148504
rect 428274 148452 428280 148504
rect 428332 148492 428338 148504
rect 522298 148492 522304 148504
rect 428332 148464 522304 148492
rect 428332 148452 428338 148464
rect 522298 148452 522304 148464
rect 522356 148452 522362 148504
rect 11698 148384 11704 148436
rect 11756 148424 11762 148436
rect 128354 148424 128360 148436
rect 11756 148396 128360 148424
rect 11756 148384 11762 148396
rect 128354 148384 128360 148396
rect 128412 148384 128418 148436
rect 133230 148384 133236 148436
rect 133288 148424 133294 148436
rect 200390 148424 200396 148436
rect 133288 148396 200396 148424
rect 133288 148384 133294 148396
rect 200390 148384 200396 148396
rect 200448 148384 200454 148436
rect 213822 148384 213828 148436
rect 213880 148424 213886 148436
rect 247770 148424 247776 148436
rect 213880 148396 247776 148424
rect 213880 148384 213886 148396
rect 247770 148384 247776 148396
rect 247828 148384 247834 148436
rect 249702 148384 249708 148436
rect 249760 148424 249766 148436
rect 268378 148424 268384 148436
rect 249760 148396 268384 148424
rect 249760 148384 249766 148396
rect 268378 148384 268384 148396
rect 268436 148384 268442 148436
rect 268930 148384 268936 148436
rect 268988 148424 268994 148436
rect 279326 148424 279332 148436
rect 268988 148396 279332 148424
rect 268988 148384 268994 148396
rect 279326 148384 279332 148396
rect 279384 148384 279390 148436
rect 286962 148384 286968 148436
rect 287020 148424 287026 148436
rect 290274 148424 290280 148436
rect 287020 148396 290280 148424
rect 287020 148384 287026 148396
rect 290274 148384 290280 148396
rect 290332 148384 290338 148436
rect 326706 148384 326712 148436
rect 326764 148424 326770 148436
rect 349246 148424 349252 148436
rect 326764 148396 349252 148424
rect 326764 148384 326770 148396
rect 349246 148384 349252 148396
rect 349304 148384 349310 148436
rect 364426 148384 364432 148436
rect 364484 148424 364490 148436
rect 413278 148424 413284 148436
rect 364484 148396 413284 148424
rect 364484 148384 364490 148396
rect 413278 148384 413284 148396
rect 413336 148384 413342 148436
rect 430298 148384 430304 148436
rect 430356 148424 430362 148436
rect 526438 148424 526444 148436
rect 430356 148396 526444 148424
rect 430356 148384 430362 148396
rect 526438 148384 526444 148396
rect 526496 148384 526502 148436
rect 7558 148316 7564 148368
rect 7616 148356 7622 148368
rect 127710 148356 127716 148368
rect 7616 148328 127716 148356
rect 7616 148316 7622 148328
rect 127710 148316 127716 148328
rect 127768 148316 127774 148368
rect 128998 148316 129004 148368
rect 129056 148356 129062 148368
rect 198366 148356 198372 148368
rect 129056 148328 198372 148356
rect 129056 148316 129062 148328
rect 198366 148316 198372 148328
rect 198424 148316 198430 148368
rect 205542 148316 205548 148368
rect 205600 148356 205606 148368
rect 242986 148356 242992 148368
rect 205600 148328 242992 148356
rect 205600 148316 205606 148328
rect 242986 148316 242992 148328
rect 243044 148316 243050 148368
rect 244918 148316 244924 148368
rect 244976 148356 244982 148368
rect 265618 148356 265624 148368
rect 244976 148328 265624 148356
rect 244976 148316 244982 148328
rect 265618 148316 265624 148328
rect 265676 148316 265682 148368
rect 267182 148316 267188 148368
rect 267240 148356 267246 148368
rect 277946 148356 277952 148368
rect 267240 148328 277952 148356
rect 267240 148316 267246 148328
rect 277946 148316 277952 148328
rect 278004 148316 278010 148368
rect 311618 148316 311624 148368
rect 311676 148356 311682 148368
rect 322198 148356 322204 148368
rect 311676 148328 322204 148356
rect 311676 148316 311682 148328
rect 322198 148316 322204 148328
rect 322256 148316 322262 148368
rect 330754 148316 330760 148368
rect 330812 148356 330818 148368
rect 356146 148356 356152 148368
rect 330812 148328 356152 148356
rect 330812 148316 330818 148328
rect 356146 148316 356152 148328
rect 356204 148316 356210 148368
rect 368566 148316 368572 148368
rect 368624 148356 368630 148368
rect 418798 148356 418804 148368
rect 368624 148328 418804 148356
rect 368624 148316 368630 148328
rect 418798 148316 418804 148328
rect 418856 148316 418862 148368
rect 426161 148359 426219 148365
rect 426161 148325 426173 148359
rect 426207 148356 426219 148359
rect 432598 148356 432604 148368
rect 426207 148328 432604 148356
rect 426207 148325 426219 148328
rect 426161 148319 426219 148325
rect 432598 148316 432604 148328
rect 432656 148316 432662 148368
rect 432690 148316 432696 148368
rect 432748 148356 432754 148368
rect 530578 148356 530584 148368
rect 432748 148328 530584 148356
rect 432748 148316 432754 148328
rect 530578 148316 530584 148328
rect 530636 148316 530642 148368
rect 111058 148248 111064 148300
rect 111116 148288 111122 148300
rect 187418 148288 187424 148300
rect 111116 148260 187424 148288
rect 111116 148248 111122 148260
rect 187418 148248 187424 148260
rect 187476 148248 187482 148300
rect 195238 148248 195244 148300
rect 195296 148288 195302 148300
rect 236086 148288 236092 148300
rect 195296 148260 236092 148288
rect 195296 148248 195302 148260
rect 236086 148248 236092 148260
rect 236144 148248 236150 148300
rect 242802 148248 242808 148300
rect 242860 148288 242866 148300
rect 264238 148288 264244 148300
rect 242860 148260 264244 148288
rect 242860 148248 242866 148260
rect 264238 148248 264244 148260
rect 264296 148248 264302 148300
rect 269022 148248 269028 148300
rect 269080 148288 269086 148300
rect 280062 148288 280068 148300
rect 269080 148260 280068 148288
rect 269080 148248 269086 148260
rect 280062 148248 280068 148260
rect 280120 148248 280126 148300
rect 402146 148248 402152 148300
rect 402204 148288 402210 148300
rect 478874 148288 478880 148300
rect 402204 148260 478880 148288
rect 402204 148248 402210 148260
rect 478874 148248 478880 148260
rect 478932 148248 478938 148300
rect 114462 148180 114468 148232
rect 114520 148220 114526 148232
rect 190178 148220 190184 148232
rect 114520 148192 190184 148220
rect 114520 148180 114526 148192
rect 190178 148180 190184 148192
rect 190236 148180 190242 148232
rect 196618 148180 196624 148232
rect 196676 148220 196682 148232
rect 225782 148220 225788 148232
rect 196676 148192 225788 148220
rect 196676 148180 196682 148192
rect 225782 148180 225788 148192
rect 225840 148180 225846 148232
rect 228358 148180 228364 148232
rect 228416 148220 228422 148232
rect 240226 148220 240232 148232
rect 228416 148192 240232 148220
rect 228416 148180 228422 148192
rect 240226 148180 240232 148192
rect 240284 148180 240290 148232
rect 246942 148180 246948 148232
rect 247000 148220 247006 148232
rect 266998 148220 267004 148232
rect 247000 148192 267004 148220
rect 247000 148180 247006 148192
rect 266998 148180 267004 148192
rect 267056 148180 267062 148232
rect 267642 148180 267648 148232
rect 267700 148220 267706 148232
rect 278682 148220 278688 148232
rect 267700 148192 278688 148220
rect 267700 148180 267706 148192
rect 278682 148180 278688 148192
rect 278740 148180 278746 148232
rect 398006 148180 398012 148232
rect 398064 148220 398070 148232
rect 471974 148220 471980 148232
rect 398064 148192 471980 148220
rect 398064 148180 398070 148192
rect 471974 148180 471980 148192
rect 472032 148180 472038 148232
rect 119430 148112 119436 148164
rect 119488 148152 119494 148164
rect 191466 148152 191472 148164
rect 119488 148124 191472 148152
rect 119488 148112 119494 148124
rect 191466 148112 191472 148124
rect 191524 148112 191530 148164
rect 197998 148112 198004 148164
rect 198056 148152 198062 148164
rect 236822 148152 236828 148164
rect 198056 148124 236828 148152
rect 198056 148112 198062 148124
rect 236822 148112 236828 148124
rect 236880 148112 236886 148164
rect 244182 148112 244188 148164
rect 244240 148152 244246 148164
rect 264606 148152 264612 148164
rect 244240 148124 264612 148152
rect 244240 148112 244246 148124
rect 264606 148112 264612 148124
rect 264664 148112 264670 148164
rect 402882 148112 402888 148164
rect 402940 148152 402946 148164
rect 475378 148152 475384 148164
rect 402940 148124 475384 148152
rect 402940 148112 402946 148124
rect 475378 148112 475384 148124
rect 475436 148112 475442 148164
rect 115198 148044 115204 148096
rect 115256 148084 115262 148096
rect 115256 148056 161474 148084
rect 115256 148044 115262 148056
rect 116578 147976 116584 148028
rect 116636 148016 116642 148028
rect 155862 148016 155868 148028
rect 116636 147988 155868 148016
rect 116636 147976 116642 147988
rect 155862 147976 155868 147988
rect 155920 147976 155926 148028
rect 122098 147908 122104 147960
rect 122156 147948 122162 147960
rect 151722 147948 151728 147960
rect 122156 147920 151728 147948
rect 122156 147908 122162 147920
rect 151722 147908 151728 147920
rect 151780 147908 151786 147960
rect 161446 147948 161474 148056
rect 170398 148044 170404 148096
rect 170456 148084 170462 148096
rect 220998 148084 221004 148096
rect 170456 148056 221004 148084
rect 170456 148044 170462 148056
rect 220998 148044 221004 148056
rect 221056 148044 221062 148096
rect 240778 148044 240784 148096
rect 240836 148084 240842 148096
rect 250530 148084 250536 148096
rect 240836 148056 250536 148084
rect 240836 148044 240842 148056
rect 250530 148044 250536 148056
rect 250588 148044 250594 148096
rect 252462 148044 252468 148096
rect 252520 148084 252526 148096
rect 269758 148084 269764 148096
rect 252520 148056 269764 148084
rect 252520 148044 252526 148056
rect 269758 148044 269764 148056
rect 269816 148044 269822 148096
rect 393958 148044 393964 148096
rect 394016 148084 394022 148096
rect 465074 148084 465080 148096
rect 394016 148056 465080 148084
rect 394016 148044 394022 148056
rect 465074 148044 465080 148056
rect 465132 148044 465138 148096
rect 162210 147976 162216 148028
rect 162268 148016 162274 148028
rect 210694 148016 210700 148028
rect 162268 147988 210700 148016
rect 162268 147976 162274 147988
rect 210694 147976 210700 147988
rect 210752 147976 210758 148028
rect 251082 147976 251088 148028
rect 251140 148016 251146 148028
rect 268654 148016 268660 148028
rect 251140 147988 268660 148016
rect 251140 147976 251146 147988
rect 268654 147976 268660 147988
rect 268712 147976 268718 148028
rect 278682 147976 278688 148028
rect 278740 148016 278746 148028
rect 285490 148016 285496 148028
rect 278740 147988 285496 148016
rect 278740 147976 278746 147988
rect 285490 147976 285496 147988
rect 285548 147976 285554 148028
rect 387058 147976 387064 148028
rect 387116 148016 387122 148028
rect 390094 148016 390100 148028
rect 387116 147988 390100 148016
rect 387116 147976 387122 147988
rect 390094 147976 390100 147988
rect 390152 147976 390158 148028
rect 401502 147976 401508 148028
rect 401560 148016 401566 148028
rect 468478 148016 468484 148028
rect 401560 147988 468484 148016
rect 401560 147976 401566 147988
rect 468478 147976 468484 147988
rect 468536 147976 468542 148028
rect 170950 147948 170956 147960
rect 161446 147920 170956 147948
rect 170950 147908 170956 147920
rect 171008 147908 171014 147960
rect 255958 147908 255964 147960
rect 256016 147948 256022 147960
rect 271414 147948 271420 147960
rect 256016 147920 271420 147948
rect 256016 147908 256022 147920
rect 271414 147908 271420 147920
rect 271472 147908 271478 147960
rect 280798 147908 280804 147960
rect 280856 147948 280862 147960
rect 286226 147948 286232 147960
rect 280856 147920 286232 147948
rect 280856 147908 280862 147920
rect 286226 147908 286232 147920
rect 286284 147908 286290 147960
rect 389818 147908 389824 147960
rect 389876 147948 389882 147960
rect 456794 147948 456800 147960
rect 389876 147920 456800 147948
rect 389876 147908 389882 147920
rect 456794 147908 456800 147920
rect 456852 147908 456858 147960
rect 150434 147840 150440 147892
rect 150492 147880 150498 147892
rect 153746 147880 153752 147892
rect 150492 147852 153752 147880
rect 150492 147840 150498 147852
rect 153746 147840 153752 147852
rect 153804 147840 153810 147892
rect 257982 147840 257988 147892
rect 258040 147880 258046 147892
rect 273162 147880 273168 147892
rect 258040 147852 273168 147880
rect 258040 147840 258046 147852
rect 273162 147840 273168 147852
rect 273220 147840 273226 147892
rect 281442 147840 281448 147892
rect 281500 147880 281506 147892
rect 286870 147880 286876 147892
rect 281500 147852 286876 147880
rect 281500 147840 281506 147852
rect 286870 147840 286876 147852
rect 286928 147840 286934 147892
rect 377490 147840 377496 147892
rect 377548 147880 377554 147892
rect 436094 147880 436100 147892
rect 377548 147852 436100 147880
rect 377548 147840 377554 147852
rect 436094 147840 436100 147852
rect 436152 147840 436158 147892
rect 208394 147772 208400 147824
rect 208452 147812 208458 147824
rect 209038 147812 209044 147824
rect 208452 147784 209044 147812
rect 208452 147772 208458 147784
rect 209038 147772 209044 147784
rect 209096 147772 209102 147824
rect 219434 147772 219440 147824
rect 219492 147812 219498 147824
rect 220078 147812 220084 147824
rect 219492 147784 220084 147812
rect 219492 147772 219498 147784
rect 220078 147772 220084 147784
rect 220136 147772 220142 147824
rect 253198 147772 253204 147824
rect 253256 147812 253262 147824
rect 266262 147812 266268 147824
rect 253256 147784 266268 147812
rect 253256 147772 253262 147784
rect 266262 147772 266268 147784
rect 266320 147772 266326 147824
rect 282822 147772 282828 147824
rect 282880 147812 282886 147824
rect 287606 147812 287612 147824
rect 282880 147784 287612 147812
rect 282880 147772 282886 147784
rect 287606 147772 287612 147784
rect 287664 147772 287670 147824
rect 289630 147812 289636 147824
rect 288268 147784 289636 147812
rect 200758 147704 200764 147756
rect 200816 147744 200822 147756
rect 204530 147744 204536 147756
rect 200816 147716 204536 147744
rect 200816 147704 200822 147716
rect 204530 147704 204536 147716
rect 204588 147704 204594 147756
rect 250438 147704 250444 147756
rect 250496 147744 250502 147756
rect 262582 147744 262588 147756
rect 250496 147716 262588 147744
rect 250496 147704 250502 147716
rect 262582 147704 262588 147716
rect 262640 147704 262646 147756
rect 285490 147704 285496 147756
rect 285548 147744 285554 147756
rect 288268 147744 288296 147784
rect 289630 147772 289636 147784
rect 289688 147772 289694 147824
rect 301958 147772 301964 147824
rect 302016 147812 302022 147824
rect 306558 147812 306564 147824
rect 302016 147784 306564 147812
rect 302016 147772 302022 147784
rect 306558 147772 306564 147784
rect 306616 147772 306622 147824
rect 308858 147772 308864 147824
rect 308916 147812 308922 147824
rect 311158 147812 311164 147824
rect 308916 147784 311164 147812
rect 308916 147772 308922 147784
rect 311158 147772 311164 147784
rect 311216 147772 311222 147824
rect 337654 147772 337660 147824
rect 337712 147812 337718 147824
rect 342898 147812 342904 147824
rect 337712 147784 342904 147812
rect 337712 147772 337718 147784
rect 342898 147772 342904 147784
rect 342956 147772 342962 147824
rect 385034 147772 385040 147824
rect 385092 147812 385098 147824
rect 429838 147812 429844 147824
rect 385092 147784 429844 147812
rect 385092 147772 385098 147784
rect 429838 147772 429844 147784
rect 429896 147772 429902 147824
rect 434438 147772 434444 147824
rect 434496 147812 434502 147824
rect 467098 147812 467104 147824
rect 434496 147784 467104 147812
rect 434496 147772 434502 147784
rect 467098 147772 467104 147784
rect 467156 147772 467162 147824
rect 285548 147716 288296 147744
rect 285548 147704 285554 147716
rect 288342 147704 288348 147756
rect 288400 147744 288406 147756
rect 291010 147744 291016 147756
rect 288400 147716 291016 147744
rect 288400 147704 288406 147716
rect 291010 147704 291016 147716
rect 291068 147704 291074 147756
rect 297818 147704 297824 147756
rect 297876 147744 297882 147756
rect 298738 147744 298744 147756
rect 297876 147716 298744 147744
rect 297876 147704 297882 147716
rect 298738 147704 298744 147716
rect 298796 147704 298802 147756
rect 301314 147704 301320 147756
rect 301372 147744 301378 147756
rect 305178 147744 305184 147756
rect 301372 147716 305184 147744
rect 301372 147704 301378 147716
rect 305178 147704 305184 147716
rect 305236 147704 305242 147756
rect 309502 147704 309508 147756
rect 309560 147744 309566 147756
rect 310422 147744 310428 147756
rect 309560 147716 310428 147744
rect 309560 147704 309566 147716
rect 310422 147704 310428 147716
rect 310480 147704 310486 147756
rect 312998 147704 313004 147756
rect 313056 147744 313062 147756
rect 313918 147744 313924 147756
rect 313056 147716 313924 147744
rect 313056 147704 313062 147716
rect 313918 147704 313924 147716
rect 313976 147704 313982 147756
rect 315022 147704 315028 147756
rect 315080 147744 315086 147756
rect 318058 147744 318064 147756
rect 315080 147716 318064 147744
rect 315080 147704 315086 147716
rect 318058 147704 318064 147716
rect 318116 147704 318122 147756
rect 332870 147704 332876 147756
rect 332928 147744 332934 147756
rect 334618 147744 334624 147756
rect 332928 147716 334624 147744
rect 332928 147704 332934 147716
rect 334618 147704 334624 147716
rect 334676 147704 334682 147756
rect 337010 147704 337016 147756
rect 337068 147744 337074 147756
rect 340138 147744 340144 147756
rect 337068 147716 340144 147744
rect 337068 147704 337074 147716
rect 340138 147704 340144 147716
rect 340196 147704 340202 147756
rect 343818 147704 343824 147756
rect 343876 147744 343882 147756
rect 345658 147744 345664 147756
rect 343876 147716 345664 147744
rect 343876 147704 343882 147716
rect 345658 147704 345664 147716
rect 345716 147704 345722 147756
rect 389174 147704 389180 147756
rect 389232 147744 389238 147756
rect 426161 147747 426219 147753
rect 426161 147744 426173 147747
rect 389232 147716 426173 147744
rect 389232 147704 389238 147716
rect 426161 147713 426173 147716
rect 426207 147713 426219 147747
rect 426161 147707 426219 147713
rect 426820 147716 430620 147744
rect 123478 147636 123484 147688
rect 123536 147676 123542 147688
rect 125594 147676 125600 147688
rect 123536 147648 125600 147676
rect 123536 147636 123542 147648
rect 125594 147636 125600 147648
rect 125652 147636 125658 147688
rect 185302 147676 185308 147688
rect 183020 147648 185308 147676
rect 106182 147568 106188 147620
rect 106240 147608 106246 147620
rect 183020 147608 183048 147648
rect 185302 147636 185308 147648
rect 185360 147636 185366 147688
rect 191098 147636 191104 147688
rect 191156 147676 191162 147688
rect 193582 147676 193588 147688
rect 191156 147648 193588 147676
rect 191156 147636 191162 147648
rect 193582 147636 193588 147648
rect 193640 147636 193646 147688
rect 202138 147636 202144 147688
rect 202196 147676 202202 147688
rect 203886 147676 203892 147688
rect 202196 147648 203892 147676
rect 202196 147636 202202 147648
rect 203886 147636 203892 147648
rect 203944 147636 203950 147688
rect 209038 147636 209044 147688
rect 209096 147676 209102 147688
rect 211430 147676 211436 147688
rect 209096 147648 211436 147676
rect 209096 147636 209102 147648
rect 211430 147636 211436 147648
rect 211488 147636 211494 147688
rect 220078 147636 220084 147688
rect 220136 147676 220142 147688
rect 221734 147676 221740 147688
rect 220136 147648 221740 147676
rect 220136 147636 220142 147648
rect 221734 147636 221740 147648
rect 221792 147636 221798 147688
rect 224218 147636 224224 147688
rect 224276 147676 224282 147688
rect 225138 147676 225144 147688
rect 224276 147648 225144 147676
rect 224276 147636 224282 147648
rect 225138 147636 225144 147648
rect 225196 147636 225202 147688
rect 232498 147636 232504 147688
rect 232556 147676 232562 147688
rect 234062 147676 234068 147688
rect 232556 147648 234068 147676
rect 232556 147636 232562 147648
rect 234062 147636 234068 147648
rect 234120 147636 234126 147688
rect 285582 147636 285588 147688
rect 285640 147676 285646 147688
rect 288986 147676 288992 147688
rect 285640 147648 288992 147676
rect 285640 147636 285646 147648
rect 288986 147636 288992 147648
rect 289044 147636 289050 147688
rect 289722 147636 289728 147688
rect 289780 147676 289786 147688
rect 291654 147676 291660 147688
rect 289780 147648 291660 147676
rect 289780 147636 289786 147648
rect 291654 147636 291660 147648
rect 291712 147636 291718 147688
rect 297174 147636 297180 147688
rect 297232 147676 297238 147688
rect 298278 147676 298284 147688
rect 297232 147648 298284 147676
rect 297232 147636 297238 147648
rect 298278 147636 298284 147648
rect 298336 147636 298342 147688
rect 298554 147636 298560 147688
rect 298612 147676 298618 147688
rect 299658 147676 299664 147688
rect 298612 147648 299664 147676
rect 298612 147636 298618 147648
rect 299658 147636 299664 147648
rect 299716 147636 299722 147688
rect 299934 147636 299940 147688
rect 299992 147676 299998 147688
rect 302418 147676 302424 147688
rect 299992 147648 302424 147676
rect 299992 147636 299998 147648
rect 302418 147636 302424 147648
rect 302476 147636 302482 147688
rect 302694 147636 302700 147688
rect 302752 147676 302758 147688
rect 303430 147676 303436 147688
rect 302752 147648 303436 147676
rect 302752 147636 302758 147648
rect 303430 147636 303436 147648
rect 303488 147636 303494 147688
rect 305454 147636 305460 147688
rect 305512 147676 305518 147688
rect 306190 147676 306196 147688
rect 305512 147648 306196 147676
rect 305512 147636 305518 147648
rect 306190 147636 306196 147648
rect 306248 147636 306254 147688
rect 306742 147636 306748 147688
rect 306800 147676 306806 147688
rect 307662 147676 307668 147688
rect 306800 147648 307668 147676
rect 306800 147636 306806 147648
rect 307662 147636 307668 147648
rect 307720 147636 307726 147688
rect 308122 147636 308128 147688
rect 308180 147676 308186 147688
rect 309778 147676 309784 147688
rect 308180 147648 309784 147676
rect 308180 147636 308186 147648
rect 309778 147636 309784 147648
rect 309836 147636 309842 147688
rect 310882 147636 310888 147688
rect 310940 147676 310946 147688
rect 311802 147676 311808 147688
rect 310940 147648 311808 147676
rect 310940 147636 310946 147648
rect 311802 147636 311808 147648
rect 311860 147636 311866 147688
rect 312262 147636 312268 147688
rect 312320 147676 312326 147688
rect 313182 147676 313188 147688
rect 312320 147648 313188 147676
rect 312320 147636 312326 147648
rect 313182 147636 313188 147648
rect 313240 147636 313246 147688
rect 313642 147636 313648 147688
rect 313700 147676 313706 147688
rect 314470 147676 314476 147688
rect 313700 147648 314476 147676
rect 313700 147636 313706 147648
rect 314470 147636 314476 147648
rect 314528 147636 314534 147688
rect 316402 147636 316408 147688
rect 316460 147676 316466 147688
rect 317230 147676 317236 147688
rect 316460 147648 317236 147676
rect 316460 147636 316466 147648
rect 317230 147636 317236 147648
rect 317288 147636 317294 147688
rect 317782 147636 317788 147688
rect 317840 147676 317846 147688
rect 318610 147676 318616 147688
rect 317840 147648 318616 147676
rect 317840 147636 317846 147648
rect 318610 147636 318616 147648
rect 318668 147636 318674 147688
rect 319162 147636 319168 147688
rect 319220 147676 319226 147688
rect 320082 147676 320088 147688
rect 319220 147648 320088 147676
rect 319220 147636 319226 147648
rect 320082 147636 320088 147648
rect 320140 147636 320146 147688
rect 320542 147636 320548 147688
rect 320600 147676 320606 147688
rect 321370 147676 321376 147688
rect 320600 147648 321376 147676
rect 320600 147636 320606 147648
rect 321370 147636 321376 147648
rect 321428 147636 321434 147688
rect 321922 147636 321928 147688
rect 321980 147676 321986 147688
rect 322842 147676 322848 147688
rect 321980 147648 322848 147676
rect 321980 147636 321986 147648
rect 322842 147636 322848 147648
rect 322900 147636 322906 147688
rect 323210 147636 323216 147688
rect 323268 147676 323274 147688
rect 324222 147676 324228 147688
rect 323268 147648 324228 147676
rect 323268 147636 323274 147648
rect 324222 147636 324228 147648
rect 324280 147636 324286 147688
rect 324590 147636 324596 147688
rect 324648 147676 324654 147688
rect 325510 147676 325516 147688
rect 324648 147648 325516 147676
rect 324648 147636 324654 147648
rect 325510 147636 325516 147648
rect 325568 147636 325574 147688
rect 325970 147636 325976 147688
rect 326028 147676 326034 147688
rect 326982 147676 326988 147688
rect 326028 147648 326988 147676
rect 326028 147636 326034 147648
rect 326982 147636 326988 147648
rect 327040 147636 327046 147688
rect 327350 147636 327356 147688
rect 327408 147676 327414 147688
rect 328270 147676 328276 147688
rect 327408 147648 328276 147676
rect 327408 147636 327414 147648
rect 328270 147636 328276 147648
rect 328328 147636 328334 147688
rect 330110 147636 330116 147688
rect 330168 147676 330174 147688
rect 331122 147676 331128 147688
rect 330168 147648 331128 147676
rect 330168 147636 330174 147648
rect 331122 147636 331128 147648
rect 331180 147636 331186 147688
rect 331490 147636 331496 147688
rect 331548 147676 331554 147688
rect 332410 147676 332416 147688
rect 331548 147648 332416 147676
rect 331548 147636 331554 147648
rect 332410 147636 332416 147648
rect 332468 147636 332474 147688
rect 334250 147636 334256 147688
rect 334308 147676 334314 147688
rect 335262 147676 335268 147688
rect 334308 147648 335268 147676
rect 334308 147636 334314 147648
rect 335262 147636 335268 147648
rect 335320 147636 335326 147688
rect 335630 147636 335636 147688
rect 335688 147676 335694 147688
rect 336550 147676 336556 147688
rect 335688 147648 336556 147676
rect 335688 147636 335694 147648
rect 336550 147636 336556 147648
rect 336608 147636 336614 147688
rect 338390 147636 338396 147688
rect 338448 147676 338454 147688
rect 339402 147676 339408 147688
rect 338448 147648 339408 147676
rect 338448 147636 338454 147648
rect 339402 147636 339408 147648
rect 339460 147636 339466 147688
rect 339678 147636 339684 147688
rect 339736 147676 339742 147688
rect 340690 147676 340696 147688
rect 339736 147648 340696 147676
rect 339736 147636 339742 147648
rect 340690 147636 340696 147648
rect 340748 147636 340754 147688
rect 341058 147636 341064 147688
rect 341116 147676 341122 147688
rect 342162 147676 342168 147688
rect 341116 147648 342168 147676
rect 341116 147636 341122 147648
rect 342162 147636 342168 147648
rect 342220 147636 342226 147688
rect 342438 147636 342444 147688
rect 342496 147676 342502 147688
rect 343542 147676 343548 147688
rect 342496 147648 343548 147676
rect 342496 147636 342502 147648
rect 343542 147636 343548 147648
rect 343600 147636 343606 147688
rect 345198 147636 345204 147688
rect 345256 147676 345262 147688
rect 346210 147676 346216 147688
rect 345256 147648 346216 147676
rect 345256 147636 345262 147648
rect 346210 147636 346216 147648
rect 346268 147636 346274 147688
rect 346578 147636 346584 147688
rect 346636 147676 346642 147688
rect 347682 147676 347688 147688
rect 346636 147648 347688 147676
rect 346636 147636 346642 147648
rect 347682 147636 347688 147648
rect 347740 147636 347746 147688
rect 350718 147636 350724 147688
rect 350776 147676 350782 147688
rect 351822 147676 351828 147688
rect 350776 147648 351828 147676
rect 350776 147636 350782 147648
rect 351822 147636 351828 147648
rect 351880 147636 351886 147688
rect 352098 147636 352104 147688
rect 352156 147676 352162 147688
rect 353202 147676 353208 147688
rect 352156 147648 353208 147676
rect 352156 147636 352162 147648
rect 353202 147636 353208 147648
rect 353260 147636 353266 147688
rect 353478 147636 353484 147688
rect 353536 147676 353542 147688
rect 354582 147676 354588 147688
rect 353536 147648 354588 147676
rect 353536 147636 353542 147648
rect 354582 147636 354588 147648
rect 354640 147636 354646 147688
rect 354858 147636 354864 147688
rect 354916 147676 354922 147688
rect 355962 147676 355968 147688
rect 354916 147648 355968 147676
rect 354916 147636 354922 147648
rect 355962 147636 355968 147648
rect 356020 147636 356026 147688
rect 357526 147636 357532 147688
rect 357584 147676 357590 147688
rect 358722 147676 358728 147688
rect 357584 147648 358728 147676
rect 357584 147636 357590 147648
rect 358722 147636 358728 147648
rect 358780 147636 358786 147688
rect 358906 147636 358912 147688
rect 358964 147676 358970 147688
rect 360102 147676 360108 147688
rect 358964 147648 360108 147676
rect 358964 147636 358970 147648
rect 360102 147636 360108 147648
rect 360160 147636 360166 147688
rect 361666 147636 361672 147688
rect 361724 147676 361730 147688
rect 362862 147676 362868 147688
rect 361724 147648 362868 147676
rect 361724 147636 361730 147648
rect 362862 147636 362868 147648
rect 362920 147636 362926 147688
rect 363046 147636 363052 147688
rect 363104 147676 363110 147688
rect 364242 147676 364248 147688
rect 363104 147648 364248 147676
rect 363104 147636 363110 147648
rect 364242 147636 364248 147648
rect 364300 147636 364306 147688
rect 365806 147636 365812 147688
rect 365864 147676 365870 147688
rect 367002 147676 367008 147688
rect 365864 147648 367008 147676
rect 365864 147636 365870 147648
rect 367002 147636 367008 147648
rect 367060 147636 367066 147688
rect 367186 147636 367192 147688
rect 367244 147676 367250 147688
rect 368382 147676 368388 147688
rect 367244 147648 368388 147676
rect 367244 147636 367250 147648
rect 368382 147636 368388 147648
rect 368440 147636 368446 147688
rect 369946 147636 369952 147688
rect 370004 147676 370010 147688
rect 371142 147676 371148 147688
rect 370004 147648 371148 147676
rect 370004 147636 370010 147648
rect 371142 147636 371148 147648
rect 371200 147636 371206 147688
rect 371326 147636 371332 147688
rect 371384 147676 371390 147688
rect 372522 147676 372528 147688
rect 371384 147648 372528 147676
rect 371384 147636 371390 147648
rect 372522 147636 372528 147648
rect 372580 147636 372586 147688
rect 373994 147636 374000 147688
rect 374052 147676 374058 147688
rect 375282 147676 375288 147688
rect 374052 147648 375288 147676
rect 374052 147636 374058 147648
rect 375282 147636 375288 147648
rect 375340 147636 375346 147688
rect 375374 147636 375380 147688
rect 375432 147676 375438 147688
rect 376662 147676 376668 147688
rect 375432 147648 376668 147676
rect 375432 147636 375438 147648
rect 376662 147636 376668 147648
rect 376720 147636 376726 147688
rect 376754 147636 376760 147688
rect 376812 147676 376818 147688
rect 378042 147676 378048 147688
rect 376812 147648 378048 147676
rect 376812 147636 376818 147648
rect 378042 147636 378048 147648
rect 378100 147636 378106 147688
rect 378134 147636 378140 147688
rect 378192 147676 378198 147688
rect 379422 147676 379428 147688
rect 378192 147648 379428 147676
rect 378192 147636 378198 147648
rect 379422 147636 379428 147648
rect 379480 147636 379486 147688
rect 379514 147636 379520 147688
rect 379572 147676 379578 147688
rect 380802 147676 380808 147688
rect 379572 147648 380808 147676
rect 379572 147636 379578 147648
rect 380802 147636 380808 147648
rect 380860 147636 380866 147688
rect 380894 147636 380900 147688
rect 380952 147676 380958 147688
rect 382090 147676 382096 147688
rect 380952 147648 382096 147676
rect 380952 147636 380958 147648
rect 382090 147636 382096 147648
rect 382148 147636 382154 147688
rect 382274 147636 382280 147688
rect 382332 147676 382338 147688
rect 383562 147676 383568 147688
rect 382332 147648 383568 147676
rect 382332 147636 382338 147648
rect 383562 147636 383568 147648
rect 383620 147636 383626 147688
rect 383654 147636 383660 147688
rect 383712 147676 383718 147688
rect 384942 147676 384948 147688
rect 383712 147648 384948 147676
rect 383712 147636 383718 147648
rect 384942 147636 384948 147648
rect 385000 147636 385006 147688
rect 386414 147636 386420 147688
rect 386472 147676 386478 147688
rect 387702 147676 387708 147688
rect 386472 147648 387708 147676
rect 386472 147636 386478 147648
rect 387702 147636 387708 147648
rect 387760 147636 387766 147688
rect 387794 147636 387800 147688
rect 387852 147676 387858 147688
rect 389082 147676 389088 147688
rect 387852 147648 389088 147676
rect 387852 147636 387858 147648
rect 389082 147636 389088 147648
rect 389140 147636 389146 147688
rect 391198 147636 391204 147688
rect 391256 147676 391262 147688
rect 392578 147676 392584 147688
rect 391256 147648 392584 147676
rect 391256 147636 391262 147648
rect 392578 147636 392584 147648
rect 392636 147636 392642 147688
rect 396626 147636 396632 147688
rect 396684 147676 396690 147688
rect 397362 147676 397368 147688
rect 396684 147648 397368 147676
rect 396684 147636 396690 147648
rect 397362 147636 397368 147648
rect 397420 147636 397426 147688
rect 400766 147636 400772 147688
rect 400824 147676 400830 147688
rect 401502 147676 401508 147688
rect 400824 147648 401508 147676
rect 400824 147636 400830 147648
rect 401502 147636 401508 147648
rect 401560 147636 401566 147688
rect 403526 147636 403532 147688
rect 403584 147676 403590 147688
rect 404262 147676 404268 147688
rect 403584 147648 404268 147676
rect 403584 147636 403590 147648
rect 404262 147636 404268 147648
rect 404320 147636 404326 147688
rect 404906 147636 404912 147688
rect 404964 147676 404970 147688
rect 404964 147648 407068 147676
rect 404964 147636 404970 147648
rect 106240 147580 183048 147608
rect 407040 147608 407068 147648
rect 411806 147636 411812 147688
rect 411864 147676 411870 147688
rect 412542 147676 412548 147688
rect 411864 147648 412548 147676
rect 411864 147636 411870 147648
rect 412542 147636 412548 147648
rect 412600 147636 412606 147688
rect 415854 147636 415860 147688
rect 415912 147676 415918 147688
rect 416590 147676 416596 147688
rect 415912 147648 416596 147676
rect 415912 147636 415918 147648
rect 416590 147636 416596 147648
rect 416648 147636 416654 147688
rect 421374 147636 421380 147688
rect 421432 147676 421438 147688
rect 422202 147676 422208 147688
rect 421432 147648 422208 147676
rect 421432 147636 421438 147648
rect 422202 147636 422208 147648
rect 422260 147636 422266 147688
rect 424134 147636 424140 147688
rect 424192 147676 424198 147688
rect 426820 147676 426848 147716
rect 424192 147648 426848 147676
rect 424192 147636 424198 147648
rect 426894 147636 426900 147688
rect 426952 147676 426958 147688
rect 427722 147676 427728 147688
rect 426952 147648 427728 147676
rect 426952 147636 426958 147648
rect 427722 147636 427728 147648
rect 427780 147636 427786 147688
rect 429562 147636 429568 147688
rect 429620 147676 429626 147688
rect 430482 147676 430488 147688
rect 429620 147648 430488 147676
rect 429620 147636 429626 147648
rect 430482 147636 430488 147648
rect 430540 147636 430546 147688
rect 430592 147676 430620 147716
rect 430942 147704 430948 147756
rect 431000 147744 431006 147756
rect 431862 147744 431868 147756
rect 431000 147716 431868 147744
rect 431000 147704 431006 147716
rect 431862 147704 431868 147716
rect 431920 147704 431926 147756
rect 433702 147704 433708 147756
rect 433760 147744 433766 147756
rect 434622 147744 434628 147756
rect 433760 147716 434628 147744
rect 433760 147704 433766 147716
rect 434622 147704 434628 147716
rect 434680 147704 434686 147756
rect 435082 147704 435088 147756
rect 435140 147744 435146 147756
rect 436002 147744 436008 147756
rect 435140 147716 436008 147744
rect 435140 147704 435146 147716
rect 436002 147704 436008 147716
rect 436060 147704 436066 147756
rect 437842 147704 437848 147756
rect 437900 147744 437906 147756
rect 438670 147744 438676 147756
rect 437900 147716 438676 147744
rect 437900 147704 437906 147716
rect 438670 147704 438676 147716
rect 438728 147704 438734 147756
rect 439222 147704 439228 147756
rect 439280 147744 439286 147756
rect 440142 147744 440148 147756
rect 439280 147716 440148 147744
rect 439280 147704 439286 147716
rect 440142 147704 440148 147716
rect 440200 147704 440206 147756
rect 441982 147704 441988 147756
rect 442040 147744 442046 147756
rect 442810 147744 442816 147756
rect 442040 147716 442816 147744
rect 442040 147704 442046 147716
rect 442810 147704 442816 147716
rect 442868 147704 442874 147756
rect 443362 147704 443368 147756
rect 443420 147744 443426 147756
rect 444282 147744 444288 147756
rect 443420 147716 444288 147744
rect 443420 147704 443426 147716
rect 444282 147704 444288 147716
rect 444340 147704 444346 147756
rect 446030 147704 446036 147756
rect 446088 147744 446094 147756
rect 447042 147744 447048 147756
rect 446088 147716 447048 147744
rect 446088 147704 446094 147716
rect 447042 147704 447048 147716
rect 447100 147704 447106 147756
rect 447410 147704 447416 147756
rect 447468 147744 447474 147756
rect 448422 147744 448428 147756
rect 447468 147716 448428 147744
rect 447468 147704 447474 147716
rect 448422 147704 448428 147716
rect 448480 147704 448486 147756
rect 450170 147704 450176 147756
rect 450228 147744 450234 147756
rect 451182 147744 451188 147756
rect 450228 147716 451188 147744
rect 450228 147704 450234 147716
rect 451182 147704 451188 147716
rect 451240 147704 451246 147756
rect 451550 147704 451556 147756
rect 451608 147744 451614 147756
rect 452562 147744 452568 147756
rect 451608 147716 452568 147744
rect 451608 147704 451614 147716
rect 452562 147704 452568 147716
rect 452620 147704 452626 147756
rect 454310 147704 454316 147756
rect 454368 147744 454374 147756
rect 455230 147744 455236 147756
rect 454368 147716 455236 147744
rect 454368 147704 454374 147716
rect 455230 147704 455236 147716
rect 455288 147704 455294 147756
rect 455690 147704 455696 147756
rect 455748 147744 455754 147756
rect 456702 147744 456708 147756
rect 455748 147716 456708 147744
rect 455748 147704 455754 147716
rect 456702 147704 456708 147716
rect 456760 147704 456766 147756
rect 458450 147704 458456 147756
rect 458508 147744 458514 147756
rect 459462 147744 459468 147756
rect 458508 147716 459468 147744
rect 458508 147704 458514 147716
rect 459462 147704 459468 147716
rect 459520 147704 459526 147756
rect 459830 147704 459836 147756
rect 459888 147744 459894 147756
rect 460842 147744 460848 147756
rect 459888 147716 460848 147744
rect 459888 147704 459894 147716
rect 460842 147704 460848 147716
rect 460900 147704 460906 147756
rect 464338 147744 464344 147756
rect 461136 147716 464344 147744
rect 461136 147676 461164 147716
rect 464338 147704 464344 147716
rect 464396 147704 464402 147756
rect 430592 147648 461164 147676
rect 461210 147636 461216 147688
rect 461268 147676 461274 147688
rect 462222 147676 462228 147688
rect 461268 147648 462228 147676
rect 461268 147636 461274 147648
rect 462222 147636 462228 147648
rect 462280 147636 462286 147688
rect 483014 147608 483020 147620
rect 407040 147580 483020 147608
rect 106240 147568 106246 147580
rect 483014 147568 483020 147580
rect 483072 147568 483078 147620
rect 99282 147500 99288 147552
rect 99340 147540 99346 147552
rect 177298 147540 177304 147552
rect 99340 147512 177304 147540
rect 99340 147500 99346 147512
rect 177298 147500 177304 147512
rect 177356 147500 177362 147552
rect 410794 147500 410800 147552
rect 410852 147540 410858 147552
rect 490006 147540 490012 147552
rect 410852 147512 490012 147540
rect 410852 147500 410858 147512
rect 490006 147500 490012 147512
rect 490064 147500 490070 147552
rect 95142 147432 95148 147484
rect 95200 147472 95206 147484
rect 178494 147472 178500 147484
rect 95200 147444 178500 147472
rect 95200 147432 95206 147444
rect 178494 147432 178500 147444
rect 178552 147432 178558 147484
rect 416682 147432 416688 147484
rect 416740 147472 416746 147484
rect 501598 147472 501604 147484
rect 416740 147444 501604 147472
rect 416740 147432 416746 147444
rect 501598 147432 501604 147444
rect 501656 147432 501662 147484
rect 88242 147364 88248 147416
rect 88300 147404 88306 147416
rect 174998 147404 175004 147416
rect 88300 147376 175004 147404
rect 88300 147364 88306 147376
rect 174998 147364 175004 147376
rect 175056 147364 175062 147416
rect 426158 147364 426164 147416
rect 426216 147404 426222 147416
rect 520274 147404 520280 147416
rect 426216 147376 520280 147404
rect 426216 147364 426222 147376
rect 520274 147364 520280 147376
rect 520332 147364 520338 147416
rect 59262 147296 59268 147348
rect 59320 147336 59326 147348
rect 154850 147336 154856 147348
rect 59320 147308 154856 147336
rect 59320 147296 59326 147308
rect 154850 147296 154856 147308
rect 154908 147296 154914 147348
rect 436462 147296 436468 147348
rect 436520 147336 436526 147348
rect 538214 147336 538220 147348
rect 436520 147308 538220 147336
rect 436520 147296 436526 147308
rect 538214 147296 538220 147308
rect 538272 147296 538278 147348
rect 62022 147228 62028 147280
rect 62080 147268 62086 147280
rect 159910 147268 159916 147280
rect 62080 147240 159916 147268
rect 62080 147228 62086 147240
rect 159910 147228 159916 147240
rect 159968 147228 159974 147280
rect 438486 147228 438492 147280
rect 438544 147268 438550 147280
rect 540238 147268 540244 147280
rect 438544 147240 540244 147268
rect 438544 147228 438550 147240
rect 540238 147228 540244 147240
rect 540296 147228 540302 147280
rect 52362 147160 52368 147212
rect 52420 147200 52426 147212
rect 150434 147200 150440 147212
rect 52420 147172 150440 147200
rect 52420 147160 52426 147172
rect 150434 147160 150440 147172
rect 150492 147160 150498 147212
rect 440602 147160 440608 147212
rect 440660 147200 440666 147212
rect 544378 147200 544384 147212
rect 440660 147172 544384 147200
rect 440660 147160 440666 147172
rect 544378 147160 544384 147172
rect 544436 147160 544442 147212
rect 43438 147092 43444 147144
rect 43496 147132 43502 147144
rect 146202 147132 146208 147144
rect 43496 147104 146208 147132
rect 43496 147092 43502 147104
rect 146202 147092 146208 147104
rect 146260 147092 146266 147144
rect 442626 147092 442632 147144
rect 442684 147132 442690 147144
rect 547874 147132 547880 147144
rect 442684 147104 547880 147132
rect 442684 147092 442690 147104
rect 547874 147092 547880 147104
rect 547932 147092 547938 147144
rect 47578 147024 47584 147076
rect 47636 147064 47642 147076
rect 150342 147064 150348 147076
rect 47636 147036 150348 147064
rect 47636 147024 47642 147036
rect 150342 147024 150348 147036
rect 150400 147024 150406 147076
rect 362954 147024 362960 147076
rect 363012 147064 363018 147076
rect 409874 147064 409880 147076
rect 363012 147036 409880 147064
rect 363012 147024 363018 147036
rect 409874 147024 409880 147036
rect 409932 147024 409938 147076
rect 444742 147024 444748 147076
rect 444800 147064 444806 147076
rect 551278 147064 551284 147076
rect 444800 147036 551284 147064
rect 444800 147024 444806 147036
rect 551278 147024 551284 147036
rect 551336 147024 551342 147076
rect 29638 146956 29644 147008
rect 29696 146996 29702 147008
rect 140038 146996 140044 147008
rect 29696 146968 140044 146996
rect 29696 146956 29702 146968
rect 140038 146956 140044 146968
rect 140096 146956 140102 147008
rect 367094 146956 367100 147008
rect 367152 146996 367158 147008
rect 416774 146996 416780 147008
rect 367152 146968 416780 146996
rect 367152 146956 367158 146968
rect 416774 146956 416780 146968
rect 416832 146956 416838 147008
rect 454954 146956 454960 147008
rect 455012 146996 455018 147008
rect 569218 146996 569224 147008
rect 455012 146968 569224 146996
rect 455012 146956 455018 146968
rect 569218 146956 569224 146968
rect 569276 146956 569282 147008
rect 21358 146888 21364 146940
rect 21416 146928 21422 146940
rect 134518 146928 134524 146940
rect 21416 146900 134524 146928
rect 21416 146888 21422 146900
rect 134518 146888 134524 146900
rect 134576 146888 134582 146940
rect 374638 146888 374644 146940
rect 374696 146928 374702 146940
rect 427814 146928 427820 146940
rect 374696 146900 427820 146928
rect 374696 146888 374702 146900
rect 427814 146888 427820 146900
rect 427872 146888 427878 146940
rect 457070 146888 457076 146940
rect 457128 146928 457134 146940
rect 572714 146928 572720 146940
rect 457128 146900 572720 146928
rect 457128 146888 457134 146900
rect 572714 146888 572720 146900
rect 572772 146888 572778 146940
rect 113082 146820 113088 146872
rect 113140 146860 113146 146872
rect 188982 146860 188988 146872
rect 113140 146832 188988 146860
rect 113140 146820 113146 146832
rect 188982 146820 188988 146832
rect 189040 146820 189046 146872
rect 179506 146276 179512 146328
rect 179564 146316 179570 146328
rect 180150 146316 180156 146328
rect 179564 146288 180156 146316
rect 179564 146276 179570 146288
rect 180150 146276 180156 146288
rect 180208 146276 180214 146328
rect 183646 146276 183652 146328
rect 183704 146316 183710 146328
rect 184382 146316 184388 146328
rect 183704 146288 184388 146316
rect 183704 146276 183710 146288
rect 184382 146276 184388 146288
rect 184440 146276 184446 146328
rect 196066 146276 196072 146328
rect 196124 146316 196130 146328
rect 196710 146316 196716 146328
rect 196124 146288 196716 146316
rect 196124 146276 196130 146288
rect 196710 146276 196716 146288
rect 196768 146276 196774 146328
rect 201494 146276 201500 146328
rect 201552 146316 201558 146328
rect 202230 146316 202236 146328
rect 201552 146288 202236 146316
rect 201552 146276 201558 146288
rect 202230 146276 202236 146288
rect 202288 146276 202294 146328
rect 216674 146276 216680 146328
rect 216732 146316 216738 146328
rect 217318 146316 217324 146328
rect 216732 146288 217324 146316
rect 216732 146276 216738 146288
rect 217318 146276 217324 146288
rect 217376 146276 217382 146328
rect 222194 146276 222200 146328
rect 222252 146316 222258 146328
rect 222838 146316 222844 146328
rect 222252 146288 222844 146316
rect 222252 146276 222258 146288
rect 222838 146276 222844 146288
rect 222896 146276 222902 146328
rect 226334 146276 226340 146328
rect 226392 146316 226398 146328
rect 226886 146316 226892 146328
rect 226392 146288 226892 146316
rect 226392 146276 226398 146288
rect 226886 146276 226892 146288
rect 226944 146276 226950 146328
rect 124122 146140 124128 146192
rect 124180 146180 124186 146192
rect 195606 146180 195612 146192
rect 124180 146152 195612 146180
rect 124180 146140 124186 146152
rect 195606 146140 195612 146152
rect 195664 146140 195670 146192
rect 76558 146072 76564 146124
rect 76616 146112 76622 146124
rect 167454 146112 167460 146124
rect 76616 146084 167460 146112
rect 76616 146072 76622 146084
rect 167454 146072 167460 146084
rect 167512 146072 167518 146124
rect 65518 146004 65524 146056
rect 65576 146044 65582 146056
rect 157242 146044 157248 146056
rect 65576 146016 157248 146044
rect 65576 146004 65582 146016
rect 157242 146004 157248 146016
rect 157300 146004 157306 146056
rect 71038 145936 71044 145988
rect 71096 145976 71102 145988
rect 163406 145976 163412 145988
rect 71096 145948 163412 145976
rect 71096 145936 71102 145948
rect 163406 145936 163412 145948
rect 163464 145936 163470 145988
rect 393222 145936 393228 145988
rect 393280 145976 393286 145988
rect 463694 145976 463700 145988
rect 393280 145948 463700 145976
rect 393280 145936 393286 145948
rect 463694 145936 463700 145948
rect 463752 145936 463758 145988
rect 50338 145868 50344 145920
rect 50396 145908 50402 145920
rect 148318 145908 148324 145920
rect 50396 145880 148324 145908
rect 50396 145868 50402 145880
rect 148318 145868 148324 145880
rect 148376 145868 148382 145920
rect 404170 145868 404176 145920
rect 404228 145908 404234 145920
rect 481634 145908 481640 145920
rect 404228 145880 481640 145908
rect 404228 145868 404234 145880
rect 481634 145868 481640 145880
rect 481692 145868 481698 145920
rect 53098 145800 53104 145852
rect 53156 145840 53162 145852
rect 153102 145840 153108 145852
rect 53156 145812 153108 145840
rect 53156 145800 53162 145812
rect 153102 145800 153108 145812
rect 153160 145800 153166 145852
rect 448790 145800 448796 145852
rect 448848 145840 448854 145852
rect 558178 145840 558184 145852
rect 448848 145812 558184 145840
rect 448848 145800 448854 145812
rect 558178 145800 558184 145812
rect 558236 145800 558242 145852
rect 39298 145732 39304 145784
rect 39356 145772 39362 145784
rect 144178 145772 144184 145784
rect 39356 145744 144184 145772
rect 39356 145732 39362 145744
rect 144178 145732 144184 145744
rect 144236 145732 144242 145784
rect 446766 145732 446772 145784
rect 446824 145772 446830 145784
rect 556246 145772 556252 145784
rect 446824 145744 556252 145772
rect 446824 145732 446830 145744
rect 556246 145732 556252 145744
rect 556304 145732 556310 145784
rect 32398 145664 32404 145716
rect 32456 145704 32462 145716
rect 137278 145704 137284 145716
rect 32456 145676 137284 145704
rect 32456 145664 32462 145676
rect 137278 145664 137284 145676
rect 137336 145664 137342 145716
rect 244274 145664 244280 145716
rect 244332 145704 244338 145716
rect 244734 145704 244740 145716
rect 244332 145676 244740 145704
rect 244332 145664 244338 145676
rect 244734 145664 244740 145676
rect 244792 145664 244798 145716
rect 450906 145664 450912 145716
rect 450964 145704 450970 145716
rect 560938 145704 560944 145716
rect 450964 145676 560944 145704
rect 450964 145664 450970 145676
rect 560938 145664 560944 145676
rect 560996 145664 561002 145716
rect 33778 145596 33784 145648
rect 33836 145636 33842 145648
rect 142062 145636 142068 145648
rect 33836 145608 142068 145636
rect 33836 145596 33842 145608
rect 142062 145596 142068 145608
rect 142120 145596 142126 145648
rect 452930 145596 452936 145648
rect 452988 145636 452994 145648
rect 565814 145636 565820 145648
rect 452988 145608 565820 145636
rect 452988 145596 452994 145608
rect 565814 145596 565820 145608
rect 565872 145596 565878 145648
rect 17218 145528 17224 145580
rect 17276 145568 17282 145580
rect 129734 145568 129740 145580
rect 17276 145540 129740 145568
rect 17276 145528 17282 145540
rect 129734 145528 129740 145540
rect 129792 145528 129798 145580
rect 390094 145528 390100 145580
rect 390152 145568 390158 145580
rect 452654 145568 452660 145580
rect 390152 145540 452660 145568
rect 390152 145528 390158 145540
rect 452654 145528 452660 145540
rect 452712 145528 452718 145580
rect 459094 145528 459100 145580
rect 459152 145568 459158 145580
rect 574738 145568 574744 145580
rect 459152 145540 574744 145568
rect 459152 145528 459158 145540
rect 574738 145528 574744 145540
rect 574796 145528 574802 145580
rect 168374 144848 168380 144900
rect 168432 144888 168438 144900
rect 169294 144888 169300 144900
rect 168432 144860 169300 144888
rect 168432 144848 168438 144860
rect 169294 144848 169300 144860
rect 169352 144848 169358 144900
rect 72418 144304 72424 144356
rect 72476 144344 72482 144356
rect 165430 144344 165436 144356
rect 72476 144316 165436 144344
rect 72476 144304 72482 144316
rect 165430 144304 165436 144316
rect 165488 144304 165494 144356
rect 68278 144236 68284 144288
rect 68336 144276 68342 144288
rect 161290 144276 161296 144288
rect 68336 144248 161296 144276
rect 68336 144236 68342 144248
rect 161290 144236 161296 144248
rect 161348 144236 161354 144288
rect 57238 144168 57244 144220
rect 57296 144208 57302 144220
rect 155126 144208 155132 144220
rect 57296 144180 155132 144208
rect 57296 144168 57302 144180
rect 155126 144168 155132 144180
rect 155184 144168 155190 144220
rect 408310 144168 408316 144220
rect 408368 144208 408374 144220
rect 489178 144208 489184 144220
rect 408368 144180 489184 144208
rect 408368 144168 408374 144180
rect 489178 144168 489184 144180
rect 489236 144168 489242 144220
rect 138014 142128 138020 142180
rect 138072 142168 138078 142180
rect 138198 142168 138204 142180
rect 138072 142140 138204 142168
rect 138072 142128 138078 142140
rect 138198 142128 138204 142140
rect 138256 142128 138262 142180
rect 140774 142128 140780 142180
rect 140832 142168 140838 142180
rect 140958 142168 140964 142180
rect 140832 142140 140964 142168
rect 140832 142128 140838 142140
rect 140958 142128 140964 142140
rect 141016 142128 141022 142180
rect 245654 142128 245660 142180
rect 245712 142168 245718 142180
rect 245838 142168 245844 142180
rect 245712 142140 245844 142168
rect 245712 142128 245718 142140
rect 245838 142128 245844 142140
rect 245896 142128 245902 142180
rect 256694 142128 256700 142180
rect 256752 142168 256758 142180
rect 256878 142168 256884 142180
rect 256752 142140 256884 142168
rect 256752 142128 256758 142140
rect 256878 142128 256884 142140
rect 256936 142128 256942 142180
rect 119982 141380 119988 141432
rect 120040 141420 120046 141432
rect 191098 141420 191104 141432
rect 120040 141392 191104 141420
rect 120040 141380 120046 141392
rect 191098 141380 191104 141392
rect 191156 141380 191162 141432
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 119338 137952 119344 137964
rect 3292 137924 119344 137952
rect 3292 137912 3298 137924
rect 119338 137912 119344 137924
rect 119396 137912 119402 137964
rect 3970 91740 3976 91792
rect 4028 91780 4034 91792
rect 123478 91780 123484 91792
rect 4028 91752 123484 91780
rect 4028 91740 4034 91752
rect 123478 91740 123484 91752
rect 123536 91740 123542 91792
rect 397270 33736 397276 33788
rect 397328 33776 397334 33788
rect 470594 33776 470600 33788
rect 397328 33748 470600 33776
rect 397328 33736 397334 33748
rect 470594 33736 470600 33748
rect 470652 33736 470658 33788
rect 471238 33056 471244 33108
rect 471296 33096 471302 33108
rect 580166 33096 580172 33108
rect 471296 33068 580172 33096
rect 471296 33056 471302 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 345658 25508 345664 25560
rect 345716 25548 345722 25560
rect 378134 25548 378140 25560
rect 345716 25520 378140 25548
rect 345716 25508 345722 25520
rect 378134 25508 378140 25520
rect 378192 25508 378198 25560
rect 161382 18572 161388 18624
rect 161440 18612 161446 18624
rect 216766 18612 216772 18624
rect 161440 18584 216772 18612
rect 161440 18572 161446 18584
rect 216766 18572 216772 18584
rect 216824 18572 216830 18624
rect 340690 18572 340696 18624
rect 340748 18612 340754 18624
rect 371234 18612 371240 18624
rect 340748 18584 371240 18612
rect 340748 18572 340754 18584
rect 371234 18572 371240 18584
rect 371292 18572 371298 18624
rect 412450 18572 412456 18624
rect 412508 18612 412514 18624
rect 496814 18612 496820 18624
rect 412508 18584 496820 18612
rect 412508 18572 412514 18584
rect 496814 18572 496820 18584
rect 496872 18572 496878 18624
rect 180702 17212 180708 17264
rect 180760 17252 180766 17264
rect 227806 17252 227812 17264
rect 180760 17224 227812 17252
rect 180760 17212 180766 17224
rect 227806 17212 227812 17224
rect 227864 17212 227870 17264
rect 383470 17212 383476 17264
rect 383528 17252 383534 17264
rect 445754 17252 445760 17264
rect 383528 17224 445760 17252
rect 383528 17212 383534 17224
rect 445754 17212 445760 17224
rect 445812 17212 445818 17264
rect 137646 15852 137652 15904
rect 137704 15892 137710 15904
rect 202138 15892 202144 15904
rect 137704 15864 202144 15892
rect 137704 15852 137710 15864
rect 202138 15852 202144 15864
rect 202196 15852 202202 15904
rect 215202 15852 215208 15904
rect 215260 15892 215266 15904
rect 248506 15892 248512 15904
rect 215260 15864 248512 15892
rect 215260 15852 215266 15864
rect 248506 15852 248512 15864
rect 248564 15852 248570 15904
rect 339310 15852 339316 15904
rect 339368 15892 339374 15904
rect 370130 15892 370136 15904
rect 339368 15864 370136 15892
rect 339368 15852 339374 15864
rect 370130 15852 370136 15864
rect 370188 15852 370194 15904
rect 395890 15852 395896 15904
rect 395948 15892 395954 15904
rect 467466 15892 467472 15904
rect 395948 15864 467472 15892
rect 395948 15852 395954 15864
rect 467466 15852 467472 15864
rect 467524 15852 467530 15904
rect 177942 14424 177948 14476
rect 178000 14464 178006 14476
rect 226426 14464 226432 14476
rect 178000 14436 226432 14464
rect 178000 14424 178006 14436
rect 226426 14424 226432 14436
rect 226484 14424 226490 14476
rect 429838 14424 429844 14476
rect 429896 14464 429902 14476
rect 448514 14464 448520 14476
rect 429896 14436 448520 14464
rect 429896 14424 429902 14436
rect 448514 14424 448520 14436
rect 448572 14424 448578 14476
rect 413278 13676 413284 13728
rect 413336 13716 413342 13728
rect 414290 13716 414296 13728
rect 413336 13688 414296 13716
rect 413336 13676 413342 13688
rect 414290 13676 414296 13688
rect 414348 13676 414354 13728
rect 151722 13064 151728 13116
rect 151780 13104 151786 13116
rect 209038 13104 209044 13116
rect 151780 13076 209044 13104
rect 151780 13064 151786 13076
rect 209038 13064 209044 13076
rect 209096 13064 209102 13116
rect 415302 13064 415308 13116
rect 415360 13104 415366 13116
rect 501322 13104 501328 13116
rect 415360 13076 501328 13104
rect 415360 13064 415366 13076
rect 501322 13064 501328 13076
rect 501380 13064 501386 13116
rect 133414 11704 133420 11756
rect 133472 11744 133478 11756
rect 200206 11744 200212 11756
rect 133472 11716 200212 11744
rect 133472 11704 133478 11716
rect 200206 11704 200212 11716
rect 200264 11704 200270 11756
rect 375190 11704 375196 11756
rect 375248 11744 375254 11756
rect 432046 11744 432052 11756
rect 375248 11716 432052 11744
rect 375248 11704 375254 11716
rect 432046 11704 432052 11716
rect 432104 11704 432110 11756
rect 54938 10276 54944 10328
rect 54996 10316 55002 10328
rect 116578 10316 116584 10328
rect 54996 10288 116584 10316
rect 54996 10276 55002 10288
rect 116578 10276 116584 10288
rect 116636 10276 116642 10328
rect 169662 10276 169668 10328
rect 169720 10316 169726 10328
rect 220078 10316 220084 10328
rect 169720 10288 220084 10316
rect 169720 10276 169726 10288
rect 220078 10276 220084 10288
rect 220136 10276 220142 10328
rect 419442 10276 419448 10328
rect 419500 10316 419506 10328
rect 508866 10316 508872 10328
rect 419500 10288 508872 10316
rect 419500 10276 419506 10288
rect 508866 10276 508872 10288
rect 508924 10276 508930 10328
rect 156598 9256 156604 9308
rect 156656 9296 156662 9308
rect 214006 9296 214012 9308
rect 156656 9268 214012 9296
rect 156656 9256 156662 9268
rect 214006 9256 214012 9268
rect 214064 9256 214070 9308
rect 153010 9188 153016 9240
rect 153068 9228 153074 9240
rect 212626 9228 212632 9240
rect 153068 9200 212632 9228
rect 153068 9188 153074 9200
rect 212626 9188 212632 9200
rect 212684 9188 212690 9240
rect 142430 9120 142436 9172
rect 142488 9160 142494 9172
rect 205726 9160 205732 9172
rect 142488 9132 205732 9160
rect 142488 9120 142494 9132
rect 205726 9120 205732 9132
rect 205784 9120 205790 9172
rect 145926 9052 145932 9104
rect 145984 9092 145990 9104
rect 208486 9092 208492 9104
rect 145984 9064 208492 9092
rect 145984 9052 145990 9064
rect 208486 9052 208492 9064
rect 208544 9052 208550 9104
rect 95050 8984 95056 9036
rect 95108 9024 95114 9036
rect 178126 9024 178132 9036
rect 95108 8996 178132 9024
rect 95108 8984 95114 8996
rect 178126 8984 178132 8996
rect 178184 8984 178190 9036
rect 60826 8916 60832 8968
rect 60884 8956 60890 8968
rect 158806 8956 158812 8968
rect 60884 8928 158812 8956
rect 60884 8916 60890 8928
rect 158806 8916 158812 8928
rect 158864 8916 158870 8968
rect 161290 8916 161296 8968
rect 161348 8956 161354 8968
rect 216674 8956 216680 8968
rect 161348 8928 216680 8956
rect 161348 8916 161354 8928
rect 216674 8916 216680 8928
rect 216732 8916 216738 8968
rect 343450 8916 343456 8968
rect 343508 8956 343514 8968
rect 377674 8956 377680 8968
rect 343508 8928 377680 8956
rect 343508 8916 343514 8928
rect 377674 8916 377680 8928
rect 377732 8916 377738 8968
rect 378042 8916 378048 8968
rect 378100 8956 378106 8968
rect 435542 8956 435548 8968
rect 378100 8928 435548 8956
rect 378100 8916 378106 8928
rect 435542 8916 435548 8928
rect 435600 8916 435606 8968
rect 116394 8236 116400 8288
rect 116452 8276 116458 8288
rect 119430 8276 119436 8288
rect 116452 8248 119436 8276
rect 116452 8236 116458 8248
rect 119430 8236 119436 8248
rect 119488 8236 119494 8288
rect 174262 8236 174268 8288
rect 174320 8276 174326 8288
rect 224218 8276 224224 8288
rect 174320 8248 224224 8276
rect 174320 8236 174326 8248
rect 224218 8236 224224 8248
rect 224276 8236 224282 8288
rect 169570 8168 169576 8220
rect 169628 8208 169634 8220
rect 222286 8208 222292 8220
rect 169628 8180 222292 8208
rect 169628 8168 169634 8180
rect 222286 8168 222292 8180
rect 222344 8168 222350 8220
rect 158898 8100 158904 8152
rect 158956 8140 158962 8152
rect 215386 8140 215392 8152
rect 158956 8112 215392 8140
rect 158956 8100 158962 8112
rect 215386 8100 215392 8112
rect 215444 8100 215450 8152
rect 147122 8032 147128 8084
rect 147180 8072 147186 8084
rect 208394 8072 208400 8084
rect 147180 8044 208400 8072
rect 147180 8032 147186 8044
rect 208394 8032 208400 8044
rect 208452 8032 208458 8084
rect 138842 7964 138848 8016
rect 138900 8004 138906 8016
rect 200758 8004 200764 8016
rect 138900 7976 200764 8004
rect 138900 7964 138906 7976
rect 200758 7964 200764 7976
rect 200816 7964 200822 8016
rect 425698 7964 425704 8016
rect 425756 8004 425762 8016
rect 439130 8004 439136 8016
rect 425756 7976 439136 8004
rect 425756 7964 425762 7976
rect 439130 7964 439136 7976
rect 439188 7964 439194 8016
rect 140038 7896 140044 7948
rect 140096 7936 140102 7948
rect 204346 7936 204352 7948
rect 140096 7908 204352 7936
rect 140096 7896 140102 7908
rect 204346 7896 204352 7908
rect 204404 7896 204410 7948
rect 414658 7896 414664 7948
rect 414716 7936 414722 7948
rect 424870 7936 424876 7948
rect 414716 7908 424876 7936
rect 414716 7896 414722 7908
rect 424870 7896 424876 7908
rect 424928 7896 424934 7948
rect 432598 7896 432604 7948
rect 432656 7936 432662 7948
rect 456886 7936 456892 7948
rect 432656 7908 456892 7936
rect 432656 7896 432662 7908
rect 456886 7896 456892 7908
rect 456944 7896 456950 7948
rect 468478 7896 468484 7948
rect 468536 7936 468542 7948
rect 478138 7936 478144 7948
rect 468536 7908 478144 7936
rect 468536 7896 468542 7908
rect 478138 7896 478144 7908
rect 478196 7896 478202 7948
rect 135254 7828 135260 7880
rect 135312 7868 135318 7880
rect 201494 7868 201500 7880
rect 135312 7840 201500 7868
rect 135312 7828 135318 7840
rect 201494 7828 201500 7840
rect 201552 7828 201558 7880
rect 382090 7828 382096 7880
rect 382148 7868 382154 7880
rect 442626 7868 442632 7880
rect 382148 7840 442632 7868
rect 382148 7828 382154 7840
rect 442626 7828 442632 7840
rect 442684 7828 442690 7880
rect 464338 7828 464344 7880
rect 464396 7868 464402 7880
rect 517146 7868 517152 7880
rect 464396 7840 517152 7868
rect 464396 7828 464402 7840
rect 517146 7828 517152 7840
rect 517204 7828 517210 7880
rect 134150 7760 134156 7812
rect 134208 7800 134214 7812
rect 201586 7800 201592 7812
rect 134208 7772 201592 7800
rect 134208 7760 134214 7772
rect 201586 7760 201592 7772
rect 201644 7760 201650 7812
rect 392578 7760 392584 7812
rect 392636 7800 392642 7812
rect 460382 7800 460388 7812
rect 392636 7772 460388 7800
rect 392636 7760 392642 7772
rect 460382 7760 460388 7772
rect 460440 7760 460446 7812
rect 467098 7760 467104 7812
rect 467156 7800 467162 7812
rect 534902 7800 534908 7812
rect 467156 7772 534908 7800
rect 467156 7760 467162 7772
rect 534902 7760 534908 7772
rect 534960 7760 534966 7812
rect 130562 7692 130568 7744
rect 130620 7732 130626 7744
rect 198826 7732 198832 7744
rect 130620 7704 198832 7732
rect 130620 7692 130626 7704
rect 198826 7692 198832 7704
rect 198884 7692 198890 7744
rect 400030 7692 400036 7744
rect 400088 7732 400094 7744
rect 474550 7732 474556 7744
rect 400088 7704 474556 7732
rect 400088 7692 400094 7704
rect 474550 7692 474556 7704
rect 474608 7692 474614 7744
rect 80882 7624 80888 7676
rect 80940 7664 80946 7676
rect 115198 7664 115204 7676
rect 80940 7636 115204 7664
rect 80940 7624 80946 7636
rect 115198 7624 115204 7636
rect 115256 7624 115262 7676
rect 126974 7624 126980 7676
rect 127032 7664 127038 7676
rect 197446 7664 197452 7676
rect 127032 7636 197452 7664
rect 127032 7624 127038 7636
rect 197446 7624 197452 7636
rect 197504 7624 197510 7676
rect 334618 7624 334624 7676
rect 334676 7664 334682 7676
rect 359918 7664 359924 7676
rect 334676 7636 359924 7664
rect 334676 7624 334682 7636
rect 359918 7624 359924 7636
rect 359976 7624 359982 7676
rect 407022 7624 407028 7676
rect 407080 7664 407086 7676
rect 487614 7664 487620 7676
rect 407080 7636 487620 7664
rect 407080 7624 407086 7636
rect 487614 7624 487620 7636
rect 487672 7624 487678 7676
rect 47854 7556 47860 7608
rect 47912 7596 47918 7608
rect 122098 7596 122104 7608
rect 47912 7568 122104 7596
rect 47912 7556 47918 7568
rect 122098 7556 122104 7568
rect 122156 7556 122162 7608
rect 125870 7556 125876 7608
rect 125928 7596 125934 7608
rect 196066 7596 196072 7608
rect 125928 7568 196072 7596
rect 125928 7556 125934 7568
rect 196066 7556 196072 7568
rect 196124 7556 196130 7608
rect 196802 7556 196808 7608
rect 196860 7596 196866 7608
rect 237466 7596 237472 7608
rect 196860 7568 237472 7596
rect 196860 7556 196866 7568
rect 237466 7556 237472 7568
rect 237524 7556 237530 7608
rect 358630 7556 358636 7608
rect 358688 7596 358694 7608
rect 403618 7596 403624 7608
rect 358688 7568 403624 7596
rect 358688 7556 358694 7568
rect 403618 7556 403624 7568
rect 403676 7556 403682 7608
rect 411162 7556 411168 7608
rect 411220 7596 411226 7608
rect 494698 7596 494704 7608
rect 411220 7568 494704 7596
rect 411220 7556 411226 7568
rect 494698 7556 494704 7568
rect 494756 7556 494762 7608
rect 129366 6876 129372 6928
rect 129424 6916 129430 6928
rect 133230 6916 133236 6928
rect 129424 6888 133236 6916
rect 129424 6876 129430 6888
rect 133230 6876 133236 6888
rect 133288 6876 133294 6928
rect 124214 6808 124220 6860
rect 124272 6848 124278 6860
rect 580166 6848 580172 6860
rect 124272 6820 580172 6848
rect 124272 6808 124278 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 97442 6740 97448 6792
rect 97500 6780 97506 6792
rect 179506 6780 179512 6792
rect 97500 6752 179512 6780
rect 97500 6740 97506 6752
rect 179506 6740 179512 6752
rect 179564 6740 179570 6792
rect 398742 6740 398748 6792
rect 398800 6780 398806 6792
rect 473446 6780 473452 6792
rect 398800 6752 473452 6780
rect 398800 6740 398806 6752
rect 473446 6740 473452 6752
rect 473504 6740 473510 6792
rect 84470 6672 84476 6724
rect 84528 6712 84534 6724
rect 172606 6712 172612 6724
rect 84528 6684 172612 6712
rect 84528 6672 84534 6684
rect 172606 6672 172612 6684
rect 172664 6672 172670 6724
rect 404262 6672 404268 6724
rect 404320 6712 404326 6724
rect 481726 6712 481732 6724
rect 404320 6684 481732 6712
rect 404320 6672 404326 6684
rect 481726 6672 481732 6684
rect 481784 6672 481790 6724
rect 77386 6604 77392 6656
rect 77444 6644 77450 6656
rect 168466 6644 168472 6656
rect 77444 6616 168472 6644
rect 77444 6604 77450 6616
rect 168466 6604 168472 6616
rect 168524 6604 168530 6656
rect 405642 6604 405648 6656
rect 405700 6644 405706 6656
rect 485222 6644 485228 6656
rect 405700 6616 485228 6644
rect 405700 6604 405706 6616
rect 485222 6604 485228 6616
rect 485280 6604 485286 6656
rect 70302 6536 70308 6588
rect 70360 6576 70366 6588
rect 164234 6576 164240 6588
rect 70360 6548 164240 6576
rect 70360 6536 70366 6548
rect 164234 6536 164240 6548
rect 164292 6536 164298 6588
rect 342070 6536 342076 6588
rect 342128 6576 342134 6588
rect 375190 6576 375196 6588
rect 342128 6548 375196 6576
rect 342128 6536 342134 6548
rect 375190 6536 375196 6548
rect 375248 6536 375254 6588
rect 408402 6536 408408 6588
rect 408460 6576 408466 6588
rect 488810 6576 488816 6588
rect 408460 6548 488816 6576
rect 408460 6536 408466 6548
rect 488810 6536 488816 6548
rect 488868 6536 488874 6588
rect 66714 6468 66720 6520
rect 66772 6508 66778 6520
rect 161566 6508 161572 6520
rect 66772 6480 161572 6508
rect 66772 6468 66778 6480
rect 161566 6468 161572 6480
rect 161624 6468 161630 6520
rect 346210 6468 346216 6520
rect 346268 6508 346274 6520
rect 381170 6508 381176 6520
rect 346268 6480 381176 6508
rect 346268 6468 346274 6480
rect 381170 6468 381176 6480
rect 381228 6468 381234 6520
rect 409782 6468 409788 6520
rect 409840 6508 409846 6520
rect 492306 6508 492312 6520
rect 409840 6480 492312 6508
rect 409840 6468 409846 6480
rect 492306 6468 492312 6480
rect 492364 6468 492370 6520
rect 63218 6400 63224 6452
rect 63276 6440 63282 6452
rect 160094 6440 160100 6452
rect 63276 6412 160100 6440
rect 63276 6400 63282 6412
rect 160094 6400 160100 6412
rect 160152 6400 160158 6452
rect 183738 6400 183744 6452
rect 183796 6440 183802 6452
rect 230566 6440 230572 6452
rect 183796 6412 230572 6440
rect 183796 6400 183802 6412
rect 230566 6400 230572 6412
rect 230624 6400 230630 6452
rect 346302 6400 346308 6452
rect 346360 6440 346366 6452
rect 382366 6440 382372 6452
rect 346360 6412 382372 6440
rect 346360 6400 346366 6412
rect 382366 6400 382372 6412
rect 382424 6400 382430 6452
rect 412542 6400 412548 6452
rect 412600 6440 412606 6452
rect 495894 6440 495900 6452
rect 412600 6412 495900 6440
rect 412600 6400 412606 6412
rect 495894 6400 495900 6412
rect 495952 6400 495958 6452
rect 59630 6332 59636 6384
rect 59688 6372 59694 6384
rect 157426 6372 157432 6384
rect 59688 6344 157432 6372
rect 59688 6332 59694 6344
rect 157426 6332 157432 6344
rect 157484 6332 157490 6384
rect 179046 6332 179052 6384
rect 179104 6372 179110 6384
rect 227714 6372 227720 6384
rect 179104 6344 227720 6372
rect 179104 6332 179110 6344
rect 227714 6332 227720 6344
rect 227772 6332 227778 6384
rect 350442 6332 350448 6384
rect 350500 6372 350506 6384
rect 389450 6372 389456 6384
rect 350500 6344 389456 6372
rect 350500 6332 350506 6344
rect 389450 6332 389456 6344
rect 389508 6332 389514 6384
rect 413922 6332 413928 6384
rect 413980 6372 413986 6384
rect 499390 6372 499396 6384
rect 413980 6344 499396 6372
rect 413980 6332 413986 6344
rect 499390 6332 499396 6344
rect 499448 6332 499454 6384
rect 56042 6264 56048 6316
rect 56100 6304 56106 6316
rect 155954 6304 155960 6316
rect 56100 6276 155960 6304
rect 56100 6264 56106 6276
rect 155954 6264 155960 6276
rect 156012 6264 156018 6316
rect 177850 6264 177856 6316
rect 177908 6304 177914 6316
rect 226334 6304 226340 6316
rect 177908 6276 226340 6304
rect 177908 6264 177914 6276
rect 226334 6264 226340 6276
rect 226392 6264 226398 6316
rect 353202 6264 353208 6316
rect 353260 6304 353266 6316
rect 393038 6304 393044 6316
rect 353260 6276 393044 6304
rect 353260 6264 353266 6276
rect 393038 6264 393044 6276
rect 393096 6264 393102 6316
rect 416590 6264 416596 6316
rect 416648 6304 416654 6316
rect 502886 6304 502892 6316
rect 416648 6276 502892 6304
rect 416648 6264 416654 6276
rect 502886 6264 502892 6276
rect 502944 6264 502950 6316
rect 52546 6196 52552 6248
rect 52604 6236 52610 6248
rect 153286 6236 153292 6248
rect 52604 6208 153292 6236
rect 52604 6196 52610 6208
rect 153286 6196 153292 6208
rect 153344 6196 153350 6248
rect 173250 6196 173256 6248
rect 173308 6236 173314 6248
rect 223666 6236 223672 6248
rect 173308 6208 223672 6236
rect 173308 6196 173314 6208
rect 223666 6196 223672 6208
rect 223724 6196 223730 6248
rect 357342 6196 357348 6248
rect 357400 6236 357406 6248
rect 400030 6236 400036 6248
rect 357400 6208 400036 6236
rect 357400 6196 357406 6208
rect 400030 6196 400036 6208
rect 400088 6196 400094 6248
rect 418062 6196 418068 6248
rect 418120 6236 418126 6248
rect 506474 6236 506480 6248
rect 418120 6208 506480 6236
rect 418120 6196 418126 6208
rect 506474 6196 506480 6208
rect 506532 6196 506538 6248
rect 48958 6128 48964 6180
rect 49016 6168 49022 6180
rect 151814 6168 151820 6180
rect 49016 6140 151820 6168
rect 49016 6128 49022 6140
rect 151814 6128 151820 6140
rect 151872 6128 151878 6180
rect 170766 6128 170772 6180
rect 170824 6168 170830 6180
rect 222194 6168 222200 6180
rect 170824 6140 222200 6168
rect 170824 6128 170830 6140
rect 222194 6128 222200 6140
rect 222252 6128 222258 6180
rect 354490 6128 354496 6180
rect 354548 6168 354554 6180
rect 396534 6168 396540 6180
rect 354548 6140 396540 6168
rect 354548 6128 354554 6140
rect 396534 6128 396540 6140
rect 396592 6128 396598 6180
rect 422110 6128 422116 6180
rect 422168 6168 422174 6180
rect 513558 6168 513564 6180
rect 422168 6140 513564 6168
rect 422168 6128 422174 6140
rect 513558 6128 513564 6140
rect 513616 6128 513622 6180
rect 101030 6060 101036 6112
rect 101088 6100 101094 6112
rect 182266 6100 182272 6112
rect 101088 6072 182272 6100
rect 101088 6060 101094 6072
rect 182266 6060 182272 6072
rect 182324 6060 182330 6112
rect 401502 6060 401508 6112
rect 401560 6100 401566 6112
rect 476942 6100 476948 6112
rect 401560 6072 476948 6100
rect 401560 6060 401566 6072
rect 476942 6060 476948 6072
rect 477000 6060 477006 6112
rect 104526 5992 104532 6044
rect 104584 6032 104590 6044
rect 183646 6032 183652 6044
rect 104584 6004 183652 6032
rect 104584 5992 104590 6004
rect 183646 5992 183652 6004
rect 183704 5992 183710 6044
rect 397362 5992 397368 6044
rect 397420 6032 397426 6044
rect 469858 6032 469864 6044
rect 397420 6004 469864 6032
rect 397420 5992 397426 6004
rect 469858 5992 469864 6004
rect 469916 5992 469922 6044
rect 108114 5924 108120 5976
rect 108172 5964 108178 5976
rect 186406 5964 186412 5976
rect 108172 5936 186412 5964
rect 108172 5924 108178 5936
rect 186406 5924 186412 5936
rect 186464 5924 186470 5976
rect 394602 5924 394608 5976
rect 394660 5964 394666 5976
rect 466270 5964 466276 5976
rect 394660 5936 466276 5964
rect 394660 5924 394666 5936
rect 466270 5924 466276 5936
rect 466328 5924 466334 5976
rect 111610 5856 111616 5908
rect 111668 5896 111674 5908
rect 187786 5896 187792 5908
rect 111668 5868 187792 5896
rect 111668 5856 111674 5868
rect 187786 5856 187792 5868
rect 187844 5856 187850 5908
rect 393222 5856 393228 5908
rect 393280 5896 393286 5908
rect 462774 5896 462780 5908
rect 393280 5868 462780 5896
rect 393280 5856 393286 5868
rect 462774 5856 462780 5868
rect 462832 5856 462838 5908
rect 115198 5788 115204 5840
rect 115256 5828 115262 5840
rect 190546 5828 190552 5840
rect 115256 5800 190552 5828
rect 115256 5788 115262 5800
rect 190546 5788 190552 5800
rect 190604 5788 190610 5840
rect 118786 5720 118792 5772
rect 118844 5760 118850 5772
rect 191926 5760 191932 5772
rect 118844 5732 191932 5760
rect 118844 5720 118850 5732
rect 191926 5720 191932 5732
rect 191984 5720 191990 5772
rect 122282 5652 122288 5704
rect 122340 5692 122346 5704
rect 194594 5692 194600 5704
rect 122340 5664 194600 5692
rect 122340 5652 122346 5664
rect 194594 5652 194600 5664
rect 194652 5652 194658 5704
rect 504358 5584 504364 5636
rect 504416 5624 504422 5636
rect 510062 5624 510068 5636
rect 504416 5596 510068 5624
rect 504416 5584 504422 5596
rect 510062 5584 510068 5596
rect 510120 5584 510126 5636
rect 91554 5516 91560 5568
rect 91612 5556 91618 5568
rect 93118 5556 93124 5568
rect 91612 5528 93124 5556
rect 91612 5516 91618 5528
rect 93118 5516 93124 5528
rect 93176 5516 93182 5568
rect 102226 5516 102232 5568
rect 102284 5556 102290 5568
rect 104158 5556 104164 5568
rect 102284 5528 104164 5556
rect 102284 5516 102290 5528
rect 104158 5516 104164 5528
rect 104216 5516 104222 5568
rect 109310 5516 109316 5568
rect 109368 5556 109374 5568
rect 111058 5556 111064 5568
rect 109368 5528 111064 5556
rect 109368 5516 109374 5528
rect 111058 5516 111064 5528
rect 111116 5516 111122 5568
rect 406378 5516 406384 5568
rect 406436 5556 406442 5568
rect 407206 5556 407212 5568
rect 406436 5528 407212 5556
rect 406436 5516 406442 5528
rect 407206 5516 407212 5528
rect 407264 5516 407270 5568
rect 475378 5516 475384 5568
rect 475436 5556 475442 5568
rect 480530 5556 480536 5568
rect 475436 5528 480536 5556
rect 475436 5516 475442 5528
rect 480530 5516 480536 5528
rect 480588 5516 480594 5568
rect 497458 5516 497464 5568
rect 497516 5556 497522 5568
rect 498194 5556 498200 5568
rect 497516 5528 498200 5556
rect 497516 5516 497522 5528
rect 498194 5516 498200 5528
rect 498252 5516 498258 5568
rect 502978 5516 502984 5568
rect 503036 5556 503042 5568
rect 505370 5556 505376 5568
rect 503036 5528 505376 5556
rect 503036 5516 503042 5528
rect 505370 5516 505376 5528
rect 505428 5516 505434 5568
rect 44266 5448 44272 5500
rect 44324 5488 44330 5500
rect 149146 5488 149152 5500
rect 44324 5460 149152 5488
rect 44324 5448 44330 5460
rect 149146 5448 149152 5460
rect 149204 5448 149210 5500
rect 189718 5448 189724 5500
rect 189776 5488 189782 5500
rect 232498 5488 232504 5500
rect 189776 5460 232504 5488
rect 189776 5448 189782 5460
rect 232498 5448 232504 5460
rect 232556 5448 232562 5500
rect 371142 5448 371148 5500
rect 371200 5488 371206 5500
rect 423766 5488 423772 5500
rect 371200 5460 423772 5488
rect 371200 5448 371206 5460
rect 423766 5448 423772 5460
rect 423824 5448 423830 5500
rect 435910 5448 435916 5500
rect 435968 5488 435974 5500
rect 537202 5488 537208 5500
rect 435968 5460 537208 5488
rect 435968 5448 435974 5460
rect 537202 5448 537208 5460
rect 537260 5448 537266 5500
rect 40678 5380 40684 5432
rect 40736 5420 40742 5432
rect 146386 5420 146392 5432
rect 40736 5392 146392 5420
rect 40736 5380 40742 5392
rect 146386 5380 146392 5392
rect 146444 5380 146450 5432
rect 186130 5380 186136 5432
rect 186188 5420 186194 5432
rect 231946 5420 231952 5432
rect 186188 5392 231952 5420
rect 186188 5380 186194 5392
rect 231946 5380 231952 5392
rect 232004 5380 232010 5432
rect 372430 5380 372436 5432
rect 372488 5420 372494 5432
rect 427262 5420 427268 5432
rect 372488 5392 427268 5420
rect 372488 5380 372494 5392
rect 427262 5380 427268 5392
rect 427320 5380 427326 5432
rect 440050 5380 440056 5432
rect 440108 5420 440114 5432
rect 544286 5420 544292 5432
rect 440108 5392 544292 5420
rect 440108 5380 440114 5392
rect 544286 5380 544292 5392
rect 544344 5380 544350 5432
rect 37182 5312 37188 5364
rect 37240 5352 37246 5364
rect 145006 5352 145012 5364
rect 37240 5324 145012 5352
rect 37240 5312 37246 5324
rect 145006 5312 145012 5324
rect 145064 5312 145070 5364
rect 166074 5312 166080 5364
rect 166132 5352 166138 5364
rect 219434 5352 219440 5364
rect 166132 5324 219440 5352
rect 166132 5312 166138 5324
rect 219434 5312 219440 5324
rect 219492 5312 219498 5364
rect 375282 5312 375288 5364
rect 375340 5352 375346 5364
rect 430850 5352 430856 5364
rect 375340 5324 430856 5352
rect 375340 5312 375346 5324
rect 430850 5312 430856 5324
rect 430908 5312 430914 5364
rect 442810 5312 442816 5364
rect 442868 5352 442874 5364
rect 547874 5352 547880 5364
rect 442868 5324 547880 5352
rect 442868 5312 442874 5324
rect 547874 5312 547880 5324
rect 547932 5312 547938 5364
rect 33594 5244 33600 5296
rect 33652 5284 33658 5296
rect 142246 5284 142252 5296
rect 33652 5256 142252 5284
rect 33652 5244 33658 5256
rect 142246 5244 142252 5256
rect 142304 5244 142310 5296
rect 164878 5244 164884 5296
rect 164936 5284 164942 5296
rect 219526 5284 219532 5296
rect 164936 5256 219532 5284
rect 164936 5244 164942 5256
rect 219526 5244 219532 5256
rect 219584 5244 219590 5296
rect 376570 5244 376576 5296
rect 376628 5284 376634 5296
rect 434438 5284 434444 5296
rect 376628 5256 434444 5284
rect 376628 5244 376634 5256
rect 434438 5244 434444 5256
rect 434496 5244 434502 5296
rect 444190 5244 444196 5296
rect 444248 5284 444254 5296
rect 551462 5284 551468 5296
rect 444248 5256 551468 5284
rect 444248 5244 444254 5256
rect 551462 5244 551468 5256
rect 551520 5244 551526 5296
rect 30098 5176 30104 5228
rect 30156 5216 30162 5228
rect 140866 5216 140872 5228
rect 30156 5188 140872 5216
rect 30156 5176 30162 5188
rect 140866 5176 140872 5188
rect 140924 5176 140930 5228
rect 149514 5176 149520 5228
rect 149572 5216 149578 5228
rect 162118 5216 162124 5228
rect 149572 5188 162124 5216
rect 149572 5176 149578 5188
rect 162118 5176 162124 5188
rect 162176 5176 162182 5228
rect 162486 5176 162492 5228
rect 162544 5216 162550 5228
rect 218146 5216 218152 5228
rect 162544 5188 218152 5216
rect 162544 5176 162550 5188
rect 218146 5176 218152 5188
rect 218204 5176 218210 5228
rect 379422 5176 379428 5228
rect 379480 5216 379486 5228
rect 437934 5216 437940 5228
rect 379480 5188 437940 5216
rect 379480 5176 379486 5188
rect 437934 5176 437940 5188
rect 437992 5176 437998 5228
rect 447042 5176 447048 5228
rect 447100 5216 447106 5228
rect 554958 5216 554964 5228
rect 447100 5188 554964 5216
rect 447100 5176 447106 5188
rect 554958 5176 554964 5188
rect 555016 5176 555022 5228
rect 26510 5108 26516 5160
rect 26568 5148 26574 5160
rect 139486 5148 139492 5160
rect 26568 5120 139492 5148
rect 26568 5108 26574 5120
rect 139486 5108 139492 5120
rect 139544 5108 139550 5160
rect 157794 5108 157800 5160
rect 157852 5148 157858 5160
rect 215294 5148 215300 5160
rect 157852 5120 215300 5148
rect 157852 5108 157858 5120
rect 215294 5108 215300 5120
rect 215352 5108 215358 5160
rect 325510 5108 325516 5160
rect 325568 5148 325574 5160
rect 345750 5148 345756 5160
rect 325568 5120 345756 5148
rect 325568 5108 325574 5120
rect 345750 5108 345756 5120
rect 345808 5108 345814 5160
rect 380710 5108 380716 5160
rect 380768 5148 380774 5160
rect 441522 5148 441528 5160
rect 380768 5120 441528 5148
rect 380768 5108 380774 5120
rect 441522 5108 441528 5120
rect 441580 5108 441586 5160
rect 448330 5108 448336 5160
rect 448388 5148 448394 5160
rect 558546 5148 558552 5160
rect 448388 5120 558552 5148
rect 448388 5108 448394 5120
rect 558546 5108 558552 5120
rect 558604 5108 558610 5160
rect 21818 5040 21824 5092
rect 21876 5080 21882 5092
rect 136634 5080 136640 5092
rect 21876 5052 136640 5080
rect 21876 5040 21882 5052
rect 136634 5040 136640 5052
rect 136692 5040 136698 5092
rect 151814 5040 151820 5092
rect 151872 5080 151878 5092
rect 211246 5080 211252 5092
rect 151872 5052 211252 5080
rect 151872 5040 151878 5052
rect 211246 5040 211252 5052
rect 211304 5040 211310 5092
rect 342898 5040 342904 5092
rect 342956 5080 342962 5092
rect 368198 5080 368204 5092
rect 342956 5052 368204 5080
rect 342956 5040 342962 5052
rect 368198 5040 368204 5052
rect 368256 5040 368262 5092
rect 383562 5040 383568 5092
rect 383620 5080 383626 5092
rect 445018 5080 445024 5092
rect 383620 5052 445024 5080
rect 383620 5040 383626 5052
rect 445018 5040 445024 5052
rect 445076 5040 445082 5092
rect 451182 5040 451188 5092
rect 451240 5080 451246 5092
rect 562042 5080 562048 5092
rect 451240 5052 562048 5080
rect 451240 5040 451246 5052
rect 562042 5040 562048 5052
rect 562100 5040 562106 5092
rect 17034 4972 17040 5024
rect 17092 5012 17098 5024
rect 17092 4984 131344 5012
rect 17092 4972 17098 4984
rect 12342 4904 12348 4956
rect 12400 4944 12406 4956
rect 131206 4944 131212 4956
rect 12400 4916 131212 4944
rect 12400 4904 12406 4916
rect 131206 4904 131212 4916
rect 131264 4904 131270 4956
rect 8754 4836 8760 4888
rect 8812 4876 8818 4888
rect 128446 4876 128452 4888
rect 8812 4848 128452 4876
rect 8812 4836 8818 4848
rect 128446 4836 128452 4848
rect 128504 4836 128510 4888
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 125686 4808 125692 4820
rect 4120 4780 125692 4808
rect 4120 4768 4126 4780
rect 125686 4768 125692 4780
rect 125744 4768 125750 4820
rect 131316 4808 131344 4984
rect 155402 4972 155408 5024
rect 155460 5012 155466 5024
rect 213914 5012 213920 5024
rect 155460 4984 213920 5012
rect 155460 4972 155466 4984
rect 213914 4972 213920 4984
rect 213972 4972 213978 5024
rect 218054 4972 218060 5024
rect 218112 5012 218118 5024
rect 240778 5012 240784 5024
rect 218112 4984 240784 5012
rect 218112 4972 218118 4984
rect 240778 4972 240784 4984
rect 240836 4972 240842 5024
rect 340138 4972 340144 5024
rect 340196 5012 340202 5024
rect 367002 5012 367008 5024
rect 340196 4984 367008 5012
rect 340196 4972 340202 4984
rect 367002 4972 367008 4984
rect 367060 4972 367066 5024
rect 387702 4972 387708 5024
rect 387760 5012 387766 5024
rect 452102 5012 452108 5024
rect 387760 4984 452108 5012
rect 387760 4972 387766 4984
rect 452102 4972 452108 4984
rect 452160 4972 452166 5024
rect 452470 4972 452476 5024
rect 452528 5012 452534 5024
rect 565630 5012 565636 5024
rect 452528 4984 565636 5012
rect 452528 4972 452534 4984
rect 565630 4972 565636 4984
rect 565688 4972 565694 5024
rect 148318 4904 148324 4956
rect 148376 4944 148382 4956
rect 209866 4944 209872 4956
rect 148376 4916 209872 4944
rect 148376 4904 148382 4916
rect 209866 4904 209872 4916
rect 209924 4904 209930 4956
rect 221550 4904 221556 4956
rect 221608 4944 221614 4956
rect 252646 4944 252652 4956
rect 221608 4916 252652 4944
rect 221608 4904 221614 4916
rect 252646 4904 252652 4916
rect 252704 4904 252710 4956
rect 336550 4904 336556 4956
rect 336608 4944 336614 4956
rect 364610 4944 364616 4956
rect 336608 4916 364616 4944
rect 336608 4904 336614 4916
rect 364610 4904 364616 4916
rect 364668 4904 364674 4956
rect 384850 4904 384856 4956
rect 384908 4944 384914 4956
rect 448606 4944 448612 4956
rect 384908 4916 448612 4944
rect 384908 4904 384914 4916
rect 448606 4904 448612 4916
rect 448664 4904 448670 4956
rect 455230 4904 455236 4956
rect 455288 4944 455294 4956
rect 569126 4944 569132 4956
rect 455288 4916 569132 4944
rect 455288 4904 455294 4916
rect 569126 4904 569132 4916
rect 569184 4904 569190 4956
rect 131758 4836 131764 4888
rect 131816 4876 131822 4888
rect 133138 4876 133144 4888
rect 131816 4848 133144 4876
rect 131816 4836 131822 4848
rect 133138 4836 133144 4848
rect 133196 4836 133202 4888
rect 136450 4836 136456 4888
rect 136508 4876 136514 4888
rect 144178 4876 144184 4888
rect 136508 4848 144184 4876
rect 136508 4836 136514 4848
rect 144178 4836 144184 4848
rect 144236 4836 144242 4888
rect 144730 4836 144736 4888
rect 144788 4876 144794 4888
rect 207106 4876 207112 4888
rect 144788 4848 207112 4876
rect 144788 4836 144794 4848
rect 207106 4836 207112 4848
rect 207164 4836 207170 4888
rect 210970 4836 210976 4888
rect 211028 4876 211034 4888
rect 245746 4876 245752 4888
rect 211028 4848 245752 4876
rect 211028 4836 211034 4848
rect 245746 4836 245752 4848
rect 245804 4836 245810 4888
rect 335170 4836 335176 4888
rect 335228 4876 335234 4888
rect 363506 4876 363512 4888
rect 335228 4848 363512 4876
rect 335228 4836 335234 4848
rect 363506 4836 363512 4848
rect 363564 4836 363570 4888
rect 377398 4836 377404 4888
rect 377456 4876 377462 4888
rect 384758 4876 384764 4888
rect 377456 4848 384764 4876
rect 377456 4836 377462 4848
rect 384758 4836 384764 4848
rect 384816 4836 384822 4888
rect 388990 4836 388996 4888
rect 389048 4876 389054 4888
rect 398193 4879 398251 4885
rect 389048 4848 398144 4876
rect 389048 4836 389054 4848
rect 133966 4808 133972 4820
rect 131316 4780 133972 4808
rect 133966 4768 133972 4780
rect 134024 4768 134030 4820
rect 141234 4768 141240 4820
rect 141292 4808 141298 4820
rect 205634 4808 205640 4820
rect 141292 4780 205640 4808
rect 141292 4768 141298 4780
rect 205634 4768 205640 4780
rect 205692 4768 205698 4820
rect 207382 4768 207388 4820
rect 207440 4808 207446 4820
rect 244366 4808 244372 4820
rect 207440 4780 244372 4808
rect 207440 4768 207446 4780
rect 244366 4768 244372 4780
rect 244424 4768 244430 4820
rect 321370 4768 321376 4820
rect 321428 4808 321434 4820
rect 338666 4808 338672 4820
rect 321428 4780 338672 4808
rect 321428 4768 321434 4780
rect 338666 4768 338672 4780
rect 338724 4768 338730 4820
rect 342162 4768 342168 4820
rect 342220 4808 342226 4820
rect 374086 4808 374092 4820
rect 342220 4780 374092 4808
rect 342220 4768 342226 4780
rect 374086 4768 374092 4780
rect 374144 4768 374150 4820
rect 390462 4768 390468 4820
rect 390520 4808 390526 4820
rect 398009 4811 398067 4817
rect 398009 4808 398021 4811
rect 390520 4780 398021 4808
rect 390520 4768 390526 4780
rect 398009 4777 398021 4780
rect 398055 4777 398067 4811
rect 398116 4808 398144 4848
rect 398193 4845 398205 4879
rect 398239 4876 398251 4879
rect 459186 4876 459192 4888
rect 398239 4848 459192 4876
rect 398239 4845 398251 4848
rect 398193 4839 398251 4845
rect 459186 4836 459192 4848
rect 459244 4836 459250 4888
rect 459462 4836 459468 4888
rect 459520 4876 459526 4888
rect 576302 4876 576308 4888
rect 459520 4848 576308 4876
rect 459520 4836 459526 4848
rect 576302 4836 576308 4848
rect 576360 4836 576366 4888
rect 455690 4808 455696 4820
rect 398116 4780 455696 4808
rect 398009 4771 398067 4777
rect 455690 4768 455696 4780
rect 455748 4768 455754 4820
rect 456610 4768 456616 4820
rect 456668 4808 456674 4820
rect 572714 4808 572720 4820
rect 456668 4780 572720 4808
rect 456668 4768 456674 4780
rect 572714 4768 572720 4780
rect 572772 4768 572778 4820
rect 65518 4700 65524 4752
rect 65576 4740 65582 4752
rect 161474 4740 161480 4752
rect 65576 4712 161480 4740
rect 65576 4700 65582 4712
rect 161474 4700 161480 4712
rect 161532 4700 161538 4752
rect 175458 4700 175464 4752
rect 175516 4740 175522 4752
rect 196618 4740 196624 4752
rect 175516 4712 196624 4740
rect 175516 4700 175522 4712
rect 196618 4700 196624 4712
rect 196676 4700 196682 4752
rect 203886 4700 203892 4752
rect 203944 4740 203950 4752
rect 241606 4740 241612 4752
rect 203944 4712 241612 4740
rect 203944 4700 203950 4712
rect 241606 4700 241612 4712
rect 241664 4700 241670 4752
rect 368290 4700 368296 4752
rect 368348 4740 368354 4752
rect 420178 4740 420184 4752
rect 368348 4712 420184 4740
rect 368348 4700 368354 4712
rect 420178 4700 420184 4712
rect 420236 4700 420242 4752
rect 438670 4700 438676 4752
rect 438728 4740 438734 4752
rect 540790 4740 540796 4752
rect 438728 4712 540796 4740
rect 438728 4700 438734 4712
rect 540790 4700 540796 4712
rect 540848 4700 540854 4752
rect 73798 4632 73804 4684
rect 73856 4672 73862 4684
rect 75178 4672 75184 4684
rect 73856 4644 75184 4672
rect 73856 4632 73862 4644
rect 75178 4632 75184 4644
rect 75236 4632 75242 4684
rect 165706 4672 165712 4684
rect 79244 4644 165712 4672
rect 72602 4564 72608 4616
rect 72660 4604 72666 4616
rect 79244 4604 79272 4644
rect 165706 4632 165712 4644
rect 165764 4632 165770 4684
rect 200298 4632 200304 4684
rect 200356 4672 200362 4684
rect 228358 4672 228364 4684
rect 200356 4644 228364 4672
rect 200356 4632 200362 4644
rect 228358 4632 228364 4644
rect 228416 4632 228422 4684
rect 364150 4632 364156 4684
rect 364208 4672 364214 4684
rect 413094 4672 413100 4684
rect 364208 4644 413100 4672
rect 364208 4632 364214 4644
rect 413094 4632 413100 4644
rect 413152 4632 413158 4684
rect 431770 4632 431776 4684
rect 431828 4672 431834 4684
rect 523773 4675 523831 4681
rect 431828 4644 523724 4672
rect 431828 4632 431834 4644
rect 162854 4604 162860 4616
rect 72660 4576 79272 4604
rect 79336 4576 162860 4604
rect 72660 4564 72666 4576
rect 69106 4496 69112 4548
rect 69164 4536 69170 4548
rect 79336 4536 79364 4576
rect 162854 4564 162860 4576
rect 162912 4564 162918 4616
rect 366910 4564 366916 4616
rect 366968 4604 366974 4616
rect 416682 4604 416688 4616
rect 366968 4576 416688 4604
rect 366968 4564 366974 4576
rect 416682 4564 416688 4576
rect 416740 4564 416746 4616
rect 434622 4564 434628 4616
rect 434680 4604 434686 4616
rect 523589 4607 523647 4613
rect 523589 4604 523601 4607
rect 434680 4576 523601 4604
rect 434680 4564 434686 4576
rect 523589 4573 523601 4576
rect 523635 4573 523647 4607
rect 523589 4567 523647 4573
rect 166994 4536 167000 4548
rect 69164 4508 79364 4536
rect 79428 4508 167000 4536
rect 69164 4496 69170 4508
rect 76190 4428 76196 4480
rect 76248 4468 76254 4480
rect 79428 4468 79456 4508
rect 166994 4496 167000 4508
rect 167052 4496 167058 4548
rect 360010 4496 360016 4548
rect 360068 4536 360074 4548
rect 406010 4536 406016 4548
rect 360068 4508 406016 4536
rect 360068 4496 360074 4508
rect 406010 4496 406016 4508
rect 406068 4496 406074 4548
rect 427630 4496 427636 4548
rect 427688 4536 427694 4548
rect 523034 4536 523040 4548
rect 427688 4508 523040 4536
rect 427688 4496 427694 4508
rect 523034 4496 523040 4508
rect 523092 4496 523098 4548
rect 523696 4536 523724 4644
rect 523773 4641 523785 4675
rect 523819 4672 523831 4675
rect 533706 4672 533712 4684
rect 523819 4644 533712 4672
rect 523819 4641 523831 4644
rect 523773 4635 523831 4641
rect 533706 4632 533712 4644
rect 533764 4632 533770 4684
rect 530118 4536 530124 4548
rect 523696 4508 530124 4536
rect 530118 4496 530124 4508
rect 530176 4496 530182 4548
rect 76248 4440 79456 4468
rect 76248 4428 76254 4440
rect 79686 4428 79692 4480
rect 79744 4468 79750 4480
rect 169846 4468 169852 4480
rect 79744 4440 169852 4468
rect 79744 4428 79750 4440
rect 169846 4428 169852 4440
rect 169904 4428 169910 4480
rect 362862 4428 362868 4480
rect 362920 4468 362926 4480
rect 409598 4468 409604 4480
rect 362920 4440 409604 4468
rect 362920 4428 362926 4440
rect 409598 4428 409604 4440
rect 409656 4428 409662 4480
rect 430482 4428 430488 4480
rect 430540 4468 430546 4480
rect 526622 4468 526628 4480
rect 430540 4440 526628 4468
rect 430540 4428 430546 4440
rect 526622 4428 526628 4440
rect 526680 4428 526686 4480
rect 83274 4360 83280 4412
rect 83332 4400 83338 4412
rect 171226 4400 171232 4412
rect 83332 4372 171232 4400
rect 83332 4360 83338 4372
rect 171226 4360 171232 4372
rect 171284 4360 171290 4412
rect 355870 4360 355876 4412
rect 355928 4400 355934 4412
rect 398926 4400 398932 4412
rect 355928 4372 398932 4400
rect 355928 4360 355934 4372
rect 398926 4360 398932 4372
rect 398984 4360 398990 4412
rect 426250 4360 426256 4412
rect 426308 4400 426314 4412
rect 519538 4400 519544 4412
rect 426308 4372 519544 4400
rect 426308 4360 426314 4372
rect 519538 4360 519544 4372
rect 519596 4360 519602 4412
rect 86862 4292 86868 4344
rect 86920 4332 86926 4344
rect 173986 4332 173992 4344
rect 86920 4304 173992 4332
rect 86920 4292 86926 4304
rect 173986 4292 173992 4304
rect 174044 4292 174050 4344
rect 358722 4292 358728 4344
rect 358780 4332 358786 4344
rect 402514 4332 402520 4344
rect 358780 4304 402520 4332
rect 358780 4292 358786 4304
rect 402514 4292 402520 4304
rect 402572 4292 402578 4344
rect 423582 4292 423588 4344
rect 423640 4332 423646 4344
rect 515950 4332 515956 4344
rect 423640 4304 515956 4332
rect 423640 4292 423646 4304
rect 515950 4292 515956 4304
rect 516008 4292 516014 4344
rect 90358 4224 90364 4276
rect 90416 4264 90422 4276
rect 175366 4264 175372 4276
rect 90416 4236 175372 4264
rect 90416 4224 90422 4236
rect 175366 4224 175372 4236
rect 175424 4224 175430 4276
rect 194410 4224 194416 4276
rect 194468 4264 194474 4276
rect 197998 4264 198004 4276
rect 194468 4236 198004 4264
rect 194468 4224 194474 4236
rect 197998 4224 198004 4236
rect 198056 4224 198062 4276
rect 354582 4224 354588 4276
rect 354640 4264 354646 4276
rect 395338 4264 395344 4276
rect 354640 4236 395344 4264
rect 354640 4224 354646 4236
rect 395338 4224 395344 4236
rect 395396 4224 395402 4276
rect 422202 4224 422208 4276
rect 422260 4264 422266 4276
rect 512454 4264 512460 4276
rect 422260 4236 512460 4264
rect 422260 4224 422266 4236
rect 512454 4224 512460 4236
rect 512512 4224 512518 4276
rect 7650 4156 7656 4208
rect 7708 4196 7714 4208
rect 11698 4196 11704 4208
rect 7708 4168 11704 4196
rect 7708 4156 7714 4168
rect 11698 4156 11704 4168
rect 11756 4156 11762 4208
rect 128170 4156 128176 4208
rect 128228 4196 128234 4208
rect 128998 4196 129004 4208
rect 128228 4168 129004 4196
rect 128228 4156 128234 4168
rect 128998 4156 129004 4168
rect 129056 4156 129062 4208
rect 143534 4156 143540 4208
rect 143592 4196 143598 4208
rect 146938 4196 146944 4208
rect 143592 4168 146944 4196
rect 143592 4156 143598 4168
rect 146938 4156 146944 4168
rect 146996 4156 147002 4208
rect 154206 4156 154212 4208
rect 154264 4196 154270 4208
rect 155218 4196 155224 4208
rect 154264 4168 155224 4196
rect 154264 4156 154270 4168
rect 155218 4156 155224 4168
rect 155276 4156 155282 4208
rect 163682 4156 163688 4208
rect 163740 4196 163746 4208
rect 166258 4196 166264 4208
rect 163740 4168 166264 4196
rect 163740 4156 163746 4168
rect 166258 4156 166264 4168
rect 166316 4156 166322 4208
rect 167178 4156 167184 4208
rect 167236 4196 167242 4208
rect 170398 4196 170404 4208
rect 167236 4168 170404 4196
rect 167236 4156 167242 4168
rect 170398 4156 170404 4168
rect 170456 4156 170462 4208
rect 171962 4156 171968 4208
rect 172020 4196 172026 4208
rect 173158 4196 173164 4208
rect 172020 4168 173164 4196
rect 172020 4156 172026 4168
rect 173158 4156 173164 4168
rect 173216 4156 173222 4208
rect 182542 4156 182548 4208
rect 182600 4196 182606 4208
rect 184198 4196 184204 4208
rect 182600 4168 184204 4196
rect 182600 4156 182606 4168
rect 184198 4156 184204 4168
rect 184256 4156 184262 4208
rect 193214 4156 193220 4208
rect 193272 4196 193278 4208
rect 195238 4196 195244 4208
rect 193272 4168 195244 4196
rect 193272 4156 193278 4168
rect 195238 4156 195244 4168
rect 195296 4156 195302 4208
rect 338758 4156 338764 4208
rect 338816 4196 338822 4208
rect 342162 4196 342168 4208
rect 338816 4168 342168 4196
rect 338816 4156 338822 4168
rect 342162 4156 342168 4168
rect 342220 4156 342226 4208
rect 389818 4156 389824 4208
rect 389876 4196 389882 4208
rect 391842 4196 391848 4208
rect 389876 4168 391848 4196
rect 389876 4156 389882 4168
rect 391842 4156 391848 4168
rect 391900 4156 391906 4208
rect 418798 4156 418804 4208
rect 418856 4196 418862 4208
rect 421374 4196 421380 4208
rect 418856 4168 421380 4196
rect 418856 4156 418862 4168
rect 421374 4156 421380 4168
rect 421432 4156 421438 4208
rect 522298 4156 522304 4208
rect 522356 4196 522362 4208
rect 524230 4196 524236 4208
rect 522356 4168 524236 4196
rect 522356 4156 522362 4168
rect 524230 4156 524236 4168
rect 524288 4156 524294 4208
rect 526438 4156 526444 4208
rect 526496 4196 526502 4208
rect 527818 4196 527824 4208
rect 526496 4168 527824 4196
rect 526496 4156 526502 4168
rect 527818 4156 527824 4168
rect 527876 4156 527882 4208
rect 530578 4156 530584 4208
rect 530636 4196 530642 4208
rect 531314 4196 531320 4208
rect 530636 4168 531320 4196
rect 530636 4156 530642 4168
rect 531314 4156 531320 4168
rect 531372 4156 531378 4208
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 18598 4128 18604 4140
rect 15988 4100 18604 4128
rect 15988 4088 15994 4100
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 45462 4088 45468 4140
rect 45520 4128 45526 4140
rect 47578 4128 47584 4140
rect 45520 4100 47584 4128
rect 45520 4088 45526 4100
rect 47578 4088 47584 4100
rect 47636 4088 47642 4140
rect 93946 4088 93952 4140
rect 94004 4128 94010 4140
rect 95142 4128 95148 4140
rect 94004 4100 95148 4128
rect 94004 4088 94010 4100
rect 95142 4088 95148 4100
rect 95200 4088 95206 4140
rect 98549 4131 98607 4137
rect 98549 4097 98561 4131
rect 98595 4128 98607 4131
rect 175274 4128 175280 4140
rect 98595 4100 175280 4128
rect 98595 4097 98607 4100
rect 98549 4091 98607 4097
rect 175274 4088 175280 4100
rect 175332 4088 175338 4140
rect 208578 4088 208584 4140
rect 208636 4128 208642 4140
rect 244274 4128 244280 4140
rect 208636 4100 244280 4128
rect 208636 4088 208642 4100
rect 244274 4088 244280 4100
rect 244332 4088 244338 4140
rect 296622 4088 296628 4140
rect 296680 4128 296686 4140
rect 297266 4128 297272 4140
rect 296680 4100 297272 4128
rect 296680 4088 296686 4100
rect 297266 4088 297272 4100
rect 297324 4088 297330 4140
rect 303522 4088 303528 4140
rect 303580 4128 303586 4140
rect 309042 4128 309048 4140
rect 303580 4100 309048 4128
rect 303580 4088 303586 4100
rect 309042 4088 309048 4100
rect 309100 4088 309106 4140
rect 315942 4088 315948 4140
rect 316000 4128 316006 4140
rect 330386 4128 330392 4140
rect 316000 4100 330392 4128
rect 316000 4088 316006 4100
rect 330386 4088 330392 4100
rect 330444 4088 330450 4140
rect 332410 4088 332416 4140
rect 332468 4128 332474 4140
rect 357526 4128 357532 4140
rect 332468 4100 357532 4128
rect 332468 4088 332474 4100
rect 357526 4088 357532 4100
rect 357584 4088 357590 4140
rect 365622 4088 365628 4140
rect 365680 4128 365686 4140
rect 415486 4128 415492 4140
rect 365680 4100 415492 4128
rect 365680 4088 365686 4100
rect 415486 4088 415492 4100
rect 415544 4088 415550 4140
rect 424778 4088 424784 4140
rect 424836 4128 424842 4140
rect 424962 4128 424968 4140
rect 424836 4100 424968 4128
rect 424836 4088 424842 4100
rect 424962 4088 424968 4100
rect 425020 4088 425026 4140
rect 437290 4088 437296 4140
rect 437348 4128 437354 4140
rect 539594 4128 539600 4140
rect 437348 4100 539600 4128
rect 437348 4088 437354 4100
rect 539594 4088 539600 4100
rect 539652 4088 539658 4140
rect 574738 4088 574744 4140
rect 574796 4128 574802 4140
rect 577406 4128 577412 4140
rect 574796 4100 577412 4128
rect 574796 4088 574802 4100
rect 577406 4088 577412 4100
rect 577464 4088 577470 4140
rect 64322 4020 64328 4072
rect 64380 4060 64386 4072
rect 68278 4060 68284 4072
rect 64380 4032 68284 4060
rect 64380 4020 64386 4032
rect 68278 4020 68284 4032
rect 68336 4020 68342 4072
rect 82078 4020 82084 4072
rect 82136 4060 82142 4072
rect 171134 4060 171140 4072
rect 82136 4032 171140 4060
rect 82136 4020 82142 4032
rect 171134 4020 171140 4032
rect 171192 4020 171198 4072
rect 206186 4020 206192 4072
rect 206244 4060 206250 4072
rect 242986 4060 242992 4072
rect 206244 4032 242992 4060
rect 206244 4020 206250 4032
rect 242986 4020 242992 4032
rect 243044 4020 243050 4072
rect 317230 4020 317236 4072
rect 317288 4060 317294 4072
rect 331582 4060 331588 4072
rect 317288 4032 331588 4060
rect 317288 4020 317294 4032
rect 331582 4020 331588 4032
rect 331640 4020 331646 4072
rect 333882 4020 333888 4072
rect 333940 4060 333946 4072
rect 361114 4060 361120 4072
rect 333940 4032 361120 4060
rect 333940 4020 333946 4032
rect 361114 4020 361120 4032
rect 361172 4020 361178 4072
rect 372522 4020 372528 4072
rect 372580 4060 372586 4072
rect 426158 4060 426164 4072
rect 372580 4032 426164 4060
rect 372580 4020 372586 4032
rect 426158 4020 426164 4032
rect 426216 4020 426222 4072
rect 440142 4020 440148 4072
rect 440200 4060 440206 4072
rect 543182 4060 543188 4072
rect 440200 4032 543188 4060
rect 440200 4020 440206 4032
rect 543182 4020 543188 4032
rect 543240 4020 543246 4072
rect 41874 3952 41880 4004
rect 41932 3992 41938 4004
rect 50338 3992 50344 4004
rect 41932 3964 50344 3992
rect 41932 3952 41938 3964
rect 50338 3952 50344 3964
rect 50396 3952 50402 4004
rect 57238 3952 57244 4004
rect 57296 3992 57302 4004
rect 65426 3992 65432 4004
rect 57296 3964 65432 3992
rect 57296 3952 57302 3964
rect 65426 3952 65432 3964
rect 65484 3952 65490 4004
rect 78582 3952 78588 4004
rect 78640 3992 78646 4004
rect 168374 3992 168380 4004
rect 78640 3964 168380 3992
rect 78640 3952 78646 3964
rect 168374 3952 168380 3964
rect 168432 3952 168438 4004
rect 201494 3952 201500 4004
rect 201552 3992 201558 4004
rect 237285 3995 237343 4001
rect 237285 3992 237297 3995
rect 201552 3964 237297 3992
rect 201552 3952 201558 3964
rect 237285 3961 237297 3964
rect 237331 3961 237343 3995
rect 241514 3992 241520 4004
rect 237285 3955 237343 3961
rect 237392 3964 241520 3992
rect 46658 3884 46664 3936
rect 46716 3924 46722 3936
rect 150526 3924 150532 3936
rect 46716 3896 150532 3924
rect 46716 3884 46722 3896
rect 150526 3884 150532 3896
rect 150584 3884 150590 3936
rect 202690 3884 202696 3936
rect 202748 3924 202754 3936
rect 237392 3924 237420 3964
rect 241514 3952 241520 3964
rect 241572 3952 241578 4004
rect 307570 3952 307576 4004
rect 307628 3992 307634 4004
rect 315209 3995 315267 4001
rect 315209 3992 315221 3995
rect 307628 3964 315221 3992
rect 307628 3952 307634 3964
rect 315209 3961 315221 3964
rect 315255 3961 315267 3995
rect 315209 3955 315267 3961
rect 318702 3952 318708 4004
rect 318760 3992 318766 4004
rect 319901 3995 319959 4001
rect 318760 3964 319852 3992
rect 318760 3952 318766 3964
rect 202748 3896 237420 3924
rect 238849 3927 238907 3933
rect 202748 3884 202754 3896
rect 238849 3893 238861 3927
rect 238895 3924 238907 3927
rect 247218 3924 247224 3936
rect 238895 3896 247224 3924
rect 238895 3893 238907 3896
rect 238849 3887 238907 3893
rect 247218 3884 247224 3896
rect 247276 3884 247282 3936
rect 310422 3884 310428 3936
rect 310480 3924 310486 3936
rect 319714 3924 319720 3936
rect 310480 3896 319720 3924
rect 310480 3884 310486 3896
rect 319714 3884 319720 3896
rect 319772 3884 319778 3936
rect 319824 3924 319852 3964
rect 319901 3961 319913 3995
rect 319947 3992 319959 3995
rect 332686 3992 332692 4004
rect 319947 3964 332692 3992
rect 319947 3961 319959 3964
rect 319901 3955 319959 3961
rect 332686 3952 332692 3964
rect 332744 3952 332750 4004
rect 335262 3952 335268 4004
rect 335320 3992 335326 4004
rect 362310 3992 362316 4004
rect 335320 3964 362316 3992
rect 335320 3952 335326 3964
rect 362310 3952 362316 3964
rect 362368 3952 362374 4004
rect 369762 3952 369768 4004
rect 369820 3992 369826 4004
rect 422570 3992 422576 4004
rect 369820 3964 422576 3992
rect 369820 3952 369826 3964
rect 422570 3952 422576 3964
rect 422628 3952 422634 4004
rect 441430 3952 441436 4004
rect 441488 3992 441494 4004
rect 546678 3992 546684 4004
rect 441488 3964 546684 3992
rect 441488 3952 441494 3964
rect 546678 3952 546684 3964
rect 546736 3952 546742 4004
rect 335078 3924 335084 3936
rect 319824 3896 335084 3924
rect 335078 3884 335084 3896
rect 335136 3884 335142 3936
rect 336642 3884 336648 3936
rect 336700 3924 336706 3936
rect 365806 3924 365812 3936
rect 336700 3896 365812 3924
rect 336700 3884 336706 3896
rect 365806 3884 365812 3896
rect 365864 3884 365870 3936
rect 373902 3884 373908 3936
rect 373960 3924 373966 3936
rect 429654 3924 429660 3936
rect 373960 3896 429660 3924
rect 373960 3884 373966 3896
rect 429654 3884 429660 3896
rect 429712 3884 429718 3936
rect 444282 3884 444288 3936
rect 444340 3924 444346 3936
rect 550266 3924 550272 3936
rect 444340 3896 550272 3924
rect 444340 3884 444346 3896
rect 550266 3884 550272 3896
rect 550324 3884 550330 3936
rect 34790 3816 34796 3868
rect 34848 3856 34854 3868
rect 39298 3856 39304 3868
rect 34848 3828 39304 3856
rect 34848 3816 34854 3828
rect 39298 3816 39304 3828
rect 39356 3816 39362 3868
rect 43070 3816 43076 3868
rect 43128 3856 43134 3868
rect 147674 3856 147680 3868
rect 43128 3828 147680 3856
rect 43128 3816 43134 3828
rect 147674 3816 147680 3828
rect 147732 3816 147738 3868
rect 199102 3816 199108 3868
rect 199160 3856 199166 3868
rect 229830 3856 229836 3868
rect 199160 3828 229836 3856
rect 199160 3816 199166 3828
rect 229830 3816 229836 3828
rect 229888 3816 229894 3868
rect 229925 3859 229983 3865
rect 229925 3825 229937 3859
rect 229971 3856 229983 3859
rect 230753 3859 230811 3865
rect 230753 3856 230765 3859
rect 229971 3828 230765 3856
rect 229971 3825 229983 3828
rect 229925 3819 229983 3825
rect 230753 3825 230765 3828
rect 230799 3825 230811 3859
rect 230753 3819 230811 3825
rect 231026 3816 231032 3868
rect 231084 3856 231090 3868
rect 231762 3856 231768 3868
rect 231084 3828 231768 3856
rect 231084 3816 231090 3828
rect 231762 3816 231768 3828
rect 231820 3816 231826 3868
rect 231857 3859 231915 3865
rect 231857 3825 231869 3859
rect 231903 3856 231915 3859
rect 237374 3856 237380 3868
rect 231903 3828 237380 3856
rect 231903 3825 231915 3828
rect 231857 3819 231915 3825
rect 237374 3816 237380 3828
rect 237432 3816 237438 3868
rect 237469 3859 237527 3865
rect 237469 3825 237481 3859
rect 237515 3856 237527 3859
rect 240226 3856 240232 3868
rect 237515 3828 240232 3856
rect 237515 3825 237527 3828
rect 237469 3819 237527 3825
rect 240226 3816 240232 3828
rect 240284 3816 240290 3868
rect 309778 3816 309784 3868
rect 309836 3856 309842 3868
rect 317322 3856 317328 3868
rect 309836 3828 317328 3856
rect 309836 3816 309842 3828
rect 317322 3816 317328 3828
rect 317380 3816 317386 3868
rect 317414 3816 317420 3868
rect 317472 3856 317478 3868
rect 319901 3859 319959 3865
rect 319901 3856 319913 3859
rect 317472 3828 319913 3856
rect 317472 3816 317478 3828
rect 319901 3825 319913 3828
rect 319947 3825 319959 3859
rect 319901 3819 319959 3825
rect 319990 3816 319996 3868
rect 320048 3856 320054 3868
rect 337470 3856 337476 3868
rect 320048 3828 337476 3856
rect 320048 3816 320054 3828
rect 337470 3816 337476 3828
rect 337528 3816 337534 3868
rect 339402 3816 339408 3868
rect 339460 3856 339466 3868
rect 369394 3856 369400 3868
rect 339460 3828 369400 3856
rect 339460 3816 339466 3828
rect 369394 3816 369400 3828
rect 369452 3816 369458 3868
rect 376662 3816 376668 3868
rect 376720 3856 376726 3868
rect 433242 3856 433248 3868
rect 376720 3828 433248 3856
rect 376720 3816 376726 3828
rect 433242 3816 433248 3828
rect 433300 3816 433306 3868
rect 445570 3816 445576 3868
rect 445628 3856 445634 3868
rect 553762 3856 553768 3868
rect 445628 3828 553768 3856
rect 445628 3816 445634 3828
rect 553762 3816 553768 3828
rect 553820 3816 553826 3868
rect 23014 3748 23020 3800
rect 23072 3788 23078 3800
rect 32398 3788 32404 3800
rect 23072 3760 32404 3788
rect 23072 3748 23078 3760
rect 32398 3748 32404 3760
rect 32456 3748 32462 3800
rect 35986 3748 35992 3800
rect 36044 3788 36050 3800
rect 143626 3788 143632 3800
rect 36044 3760 143632 3788
rect 36044 3748 36050 3760
rect 143626 3748 143632 3760
rect 143684 3748 143690 3800
rect 197906 3748 197912 3800
rect 197964 3788 197970 3800
rect 229741 3791 229799 3797
rect 229741 3788 229753 3791
rect 197964 3760 229753 3788
rect 197964 3748 197970 3760
rect 229741 3757 229753 3760
rect 229787 3757 229799 3791
rect 229741 3751 229799 3757
rect 230017 3791 230075 3797
rect 230017 3757 230029 3791
rect 230063 3788 230075 3791
rect 238754 3788 238760 3800
rect 230063 3760 238760 3788
rect 230063 3757 230075 3760
rect 230017 3751 230075 3757
rect 238754 3748 238760 3760
rect 238812 3748 238818 3800
rect 245194 3748 245200 3800
rect 245252 3788 245258 3800
rect 253198 3788 253204 3800
rect 245252 3760 253204 3788
rect 245252 3748 245258 3760
rect 253198 3748 253204 3760
rect 253256 3748 253262 3800
rect 283098 3748 283104 3800
rect 283156 3788 283162 3800
rect 287146 3788 287152 3800
rect 283156 3760 287152 3788
rect 283156 3748 283162 3760
rect 287146 3748 287152 3760
rect 287204 3748 287210 3800
rect 304810 3748 304816 3800
rect 304868 3788 304874 3800
rect 310238 3788 310244 3800
rect 304868 3760 310244 3788
rect 304868 3748 304874 3760
rect 310238 3748 310244 3760
rect 310296 3748 310302 3800
rect 311802 3748 311808 3800
rect 311860 3788 311866 3800
rect 322106 3788 322112 3800
rect 311860 3760 322112 3788
rect 311860 3748 311866 3760
rect 322106 3748 322112 3760
rect 322164 3748 322170 3800
rect 322842 3748 322848 3800
rect 322900 3788 322906 3800
rect 340966 3788 340972 3800
rect 322900 3760 340972 3788
rect 322900 3748 322906 3760
rect 340966 3748 340972 3760
rect 341024 3748 341030 3800
rect 343542 3748 343548 3800
rect 343600 3788 343606 3800
rect 376478 3788 376484 3800
rect 343600 3760 376484 3788
rect 343600 3748 343606 3760
rect 376478 3748 376484 3760
rect 376536 3748 376542 3800
rect 380802 3748 380808 3800
rect 380860 3788 380866 3800
rect 440326 3788 440332 3800
rect 380860 3760 440332 3788
rect 380860 3748 380866 3760
rect 440326 3748 440332 3760
rect 440384 3748 440390 3800
rect 448422 3748 448428 3800
rect 448480 3788 448486 3800
rect 557350 3788 557356 3800
rect 448480 3760 557356 3788
rect 448480 3748 448486 3760
rect 557350 3748 557356 3760
rect 557408 3748 557414 3800
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 35158 3720 35164 3732
rect 19484 3692 35164 3720
rect 19484 3680 19490 3692
rect 35158 3680 35164 3692
rect 35216 3680 35222 3732
rect 39574 3680 39580 3732
rect 39632 3720 39638 3732
rect 146294 3720 146300 3732
rect 39632 3692 146300 3720
rect 39632 3680 39638 3692
rect 146294 3680 146300 3692
rect 146352 3680 146358 3732
rect 192018 3680 192024 3732
rect 192076 3720 192082 3732
rect 192076 3692 229784 3720
rect 192076 3680 192082 3692
rect 32398 3612 32404 3664
rect 32456 3652 32462 3664
rect 142154 3652 142160 3664
rect 32456 3624 142160 3652
rect 32456 3612 32462 3624
rect 142154 3612 142160 3624
rect 142212 3612 142218 3664
rect 195606 3612 195612 3664
rect 195664 3652 195670 3664
rect 226518 3652 226524 3664
rect 195664 3624 226524 3652
rect 195664 3612 195670 3624
rect 226518 3612 226524 3624
rect 226576 3612 226582 3664
rect 226613 3655 226671 3661
rect 226613 3621 226625 3655
rect 226659 3652 226671 3655
rect 229649 3655 229707 3661
rect 229649 3652 229661 3655
rect 226659 3624 229661 3652
rect 226659 3621 226671 3624
rect 226613 3615 226671 3621
rect 229649 3621 229661 3624
rect 229695 3621 229707 3655
rect 229649 3615 229707 3621
rect 566 3544 572 3596
rect 624 3584 630 3596
rect 14458 3584 14464 3596
rect 624 3556 14464 3584
rect 624 3544 630 3556
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 25498 3584 25504 3596
rect 16546 3556 25504 3584
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3970 3516 3976 3528
rect 2924 3488 3976 3516
rect 2924 3476 2930 3488
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 16546 3516 16574 3556
rect 25498 3544 25504 3556
rect 25556 3544 25562 3596
rect 28902 3544 28908 3596
rect 28960 3584 28966 3596
rect 140958 3584 140964 3596
rect 28960 3556 140964 3584
rect 28960 3544 28966 3556
rect 140958 3544 140964 3556
rect 141016 3544 141022 3596
rect 188522 3544 188528 3596
rect 188580 3584 188586 3596
rect 226337 3587 226395 3593
rect 226337 3584 226349 3587
rect 188580 3556 226349 3584
rect 188580 3544 188586 3556
rect 226337 3553 226349 3556
rect 226383 3553 226395 3587
rect 229756 3584 229784 3692
rect 229922 3680 229928 3732
rect 229980 3720 229986 3732
rect 238846 3720 238852 3732
rect 229980 3692 238852 3720
rect 229980 3680 229986 3692
rect 238846 3680 238852 3692
rect 238904 3680 238910 3732
rect 239306 3680 239312 3732
rect 239364 3720 239370 3732
rect 250438 3720 250444 3732
rect 239364 3692 250444 3720
rect 239364 3680 239370 3692
rect 250438 3680 250444 3692
rect 250496 3680 250502 3732
rect 252370 3680 252376 3732
rect 252428 3720 252434 3732
rect 269206 3720 269212 3732
rect 252428 3692 269212 3720
rect 252428 3680 252434 3692
rect 269206 3680 269212 3692
rect 269264 3680 269270 3732
rect 310330 3680 310336 3732
rect 310388 3720 310394 3732
rect 315117 3723 315175 3729
rect 315117 3720 315129 3723
rect 310388 3692 315129 3720
rect 310388 3680 310394 3692
rect 315117 3689 315129 3692
rect 315163 3689 315175 3723
rect 315117 3683 315175 3689
rect 315209 3723 315267 3729
rect 315209 3689 315221 3723
rect 315255 3720 315267 3723
rect 316218 3720 316224 3732
rect 315255 3692 316224 3720
rect 315255 3689 315267 3692
rect 315209 3683 315267 3689
rect 316218 3680 316224 3692
rect 316276 3680 316282 3732
rect 321462 3680 321468 3732
rect 321520 3720 321526 3732
rect 339862 3720 339868 3732
rect 321520 3692 339868 3720
rect 321520 3680 321526 3692
rect 339862 3680 339868 3692
rect 339920 3680 339926 3732
rect 340782 3680 340788 3732
rect 340840 3720 340846 3732
rect 372890 3720 372896 3732
rect 340840 3692 372896 3720
rect 340840 3680 340846 3692
rect 372890 3680 372896 3692
rect 372948 3680 372954 3732
rect 382182 3680 382188 3732
rect 382240 3720 382246 3732
rect 443822 3720 443828 3732
rect 382240 3692 443828 3720
rect 382240 3680 382246 3692
rect 443822 3680 443828 3692
rect 443880 3680 443886 3732
rect 449710 3680 449716 3732
rect 449768 3720 449774 3732
rect 560846 3720 560852 3732
rect 449768 3692 560852 3720
rect 449768 3680 449774 3692
rect 560846 3680 560852 3692
rect 560904 3680 560910 3732
rect 229830 3612 229836 3664
rect 229888 3652 229894 3664
rect 236089 3655 236147 3661
rect 236089 3652 236101 3655
rect 229888 3624 236101 3652
rect 229888 3612 229894 3624
rect 236089 3621 236101 3624
rect 236135 3621 236147 3655
rect 236089 3615 236147 3621
rect 238110 3612 238116 3664
rect 238168 3652 238174 3664
rect 238662 3652 238668 3664
rect 238168 3624 238668 3652
rect 238168 3612 238174 3624
rect 238662 3612 238668 3624
rect 238720 3612 238726 3664
rect 238757 3655 238815 3661
rect 238757 3621 238769 3655
rect 238803 3652 238815 3655
rect 245838 3652 245844 3664
rect 238803 3624 245844 3652
rect 238803 3621 238815 3624
rect 238757 3615 238815 3621
rect 245838 3612 245844 3624
rect 245896 3612 245902 3664
rect 247586 3612 247592 3664
rect 247644 3652 247650 3664
rect 266446 3652 266452 3664
rect 247644 3624 266452 3652
rect 247644 3612 247650 3624
rect 266446 3612 266452 3624
rect 266504 3612 266510 3664
rect 304902 3612 304908 3664
rect 304960 3652 304966 3664
rect 311434 3652 311440 3664
rect 304960 3624 311440 3652
rect 304960 3612 304966 3624
rect 311434 3612 311440 3624
rect 311492 3612 311498 3664
rect 313182 3612 313188 3664
rect 313240 3652 313246 3664
rect 324406 3652 324412 3664
rect 313240 3624 324412 3652
rect 313240 3612 313246 3624
rect 324406 3612 324412 3624
rect 324464 3612 324470 3664
rect 325602 3612 325608 3664
rect 325660 3652 325666 3664
rect 346946 3652 346952 3664
rect 325660 3624 346952 3652
rect 325660 3612 325666 3624
rect 346946 3612 346952 3624
rect 347004 3612 347010 3664
rect 347682 3612 347688 3664
rect 347740 3652 347746 3664
rect 383562 3652 383568 3664
rect 347740 3624 383568 3652
rect 347740 3612 347746 3624
rect 383562 3612 383568 3624
rect 383620 3612 383626 3664
rect 384942 3612 384948 3664
rect 385000 3652 385006 3664
rect 447410 3652 447416 3664
rect 385000 3624 447416 3652
rect 385000 3612 385006 3624
rect 447410 3612 447416 3624
rect 447468 3612 447474 3664
rect 452562 3612 452568 3664
rect 452620 3652 452626 3664
rect 564434 3652 564440 3664
rect 452620 3624 564440 3652
rect 452620 3612 452626 3624
rect 564434 3612 564440 3624
rect 564492 3612 564498 3664
rect 234706 3584 234712 3596
rect 226337 3547 226395 3553
rect 226444 3556 229416 3584
rect 229756 3556 234712 3584
rect 13596 3488 16574 3516
rect 13596 3476 13602 3488
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 21358 3516 21364 3528
rect 18288 3488 21364 3516
rect 18288 3476 18294 3488
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 138106 3516 138112 3528
rect 25372 3488 138112 3516
rect 25372 3476 25378 3488
rect 138106 3476 138112 3488
rect 138164 3476 138170 3528
rect 150618 3476 150624 3528
rect 150676 3516 150682 3528
rect 151722 3516 151728 3528
rect 150676 3488 151728 3516
rect 150676 3476 150682 3488
rect 151722 3476 151728 3488
rect 151780 3476 151786 3528
rect 160094 3476 160100 3528
rect 160152 3516 160158 3528
rect 161382 3516 161388 3528
rect 160152 3488 161388 3516
rect 160152 3476 160158 3488
rect 161382 3476 161388 3488
rect 161440 3476 161446 3528
rect 168374 3476 168380 3528
rect 168432 3516 168438 3528
rect 169662 3516 169668 3528
rect 168432 3488 169668 3516
rect 168432 3476 168438 3488
rect 169662 3476 169668 3488
rect 169720 3476 169726 3528
rect 176654 3476 176660 3528
rect 176712 3516 176718 3528
rect 177942 3516 177948 3528
rect 176712 3488 177948 3516
rect 176712 3476 176718 3488
rect 177942 3476 177948 3488
rect 178000 3476 178006 3528
rect 180242 3476 180248 3528
rect 180300 3516 180306 3528
rect 180702 3516 180708 3528
rect 180300 3488 180708 3516
rect 180300 3476 180306 3488
rect 180702 3476 180708 3488
rect 180760 3476 180766 3528
rect 184934 3476 184940 3528
rect 184992 3516 184998 3528
rect 226444 3516 226472 3556
rect 184992 3488 226472 3516
rect 184992 3476 184998 3488
rect 226518 3476 226524 3528
rect 226576 3516 226582 3528
rect 229189 3519 229247 3525
rect 229189 3516 229201 3519
rect 226576 3488 229201 3516
rect 226576 3476 226582 3488
rect 229189 3485 229201 3488
rect 229235 3485 229247 3519
rect 229189 3479 229247 3485
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 22738 3448 22744 3460
rect 1728 3420 22744 3448
rect 1728 3408 1734 3420
rect 22738 3408 22744 3420
rect 22796 3408 22802 3460
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 138198 3448 138204 3460
rect 24268 3420 138204 3448
rect 24268 3408 24274 3420
rect 138198 3408 138204 3420
rect 138256 3408 138262 3460
rect 181438 3408 181444 3460
rect 181496 3448 181502 3460
rect 229278 3448 229284 3460
rect 181496 3420 229284 3448
rect 181496 3408 181502 3420
rect 229278 3408 229284 3420
rect 229336 3408 229342 3460
rect 229388 3448 229416 3556
rect 234706 3544 234712 3556
rect 234764 3544 234770 3596
rect 235810 3544 235816 3596
rect 235868 3584 235874 3596
rect 260926 3584 260932 3596
rect 235868 3556 260932 3584
rect 235868 3544 235874 3556
rect 260926 3544 260932 3556
rect 260984 3544 260990 3596
rect 267734 3544 267740 3596
rect 267792 3584 267798 3596
rect 268930 3584 268936 3596
rect 267792 3556 268936 3584
rect 267792 3544 267798 3556
rect 268930 3544 268936 3556
rect 268988 3544 268994 3596
rect 276014 3544 276020 3596
rect 276072 3584 276078 3596
rect 277210 3584 277216 3596
rect 276072 3556 277216 3584
rect 276072 3544 276078 3556
rect 277210 3544 277216 3556
rect 277268 3544 277274 3596
rect 306190 3544 306196 3596
rect 306248 3584 306254 3596
rect 312630 3584 312636 3596
rect 306248 3556 312636 3584
rect 306248 3544 306254 3556
rect 312630 3544 312636 3556
rect 312688 3544 312694 3596
rect 314562 3544 314568 3596
rect 314620 3584 314626 3596
rect 327994 3584 328000 3596
rect 314620 3556 328000 3584
rect 314620 3544 314626 3556
rect 327994 3544 328000 3556
rect 328052 3544 328058 3596
rect 328362 3544 328368 3596
rect 328420 3584 328426 3596
rect 351638 3584 351644 3596
rect 328420 3556 351644 3584
rect 328420 3544 328426 3556
rect 351638 3544 351644 3556
rect 351696 3544 351702 3596
rect 351822 3544 351828 3596
rect 351880 3584 351886 3596
rect 390646 3584 390652 3596
rect 351880 3556 390652 3584
rect 351880 3544 351886 3556
rect 390646 3544 390652 3556
rect 390704 3544 390710 3596
rect 391750 3544 391756 3596
rect 391808 3584 391814 3596
rect 461578 3584 461584 3596
rect 391808 3556 461584 3584
rect 391808 3544 391814 3556
rect 461578 3544 461584 3556
rect 461636 3544 461642 3596
rect 462222 3544 462228 3596
rect 462280 3584 462286 3596
rect 582190 3584 582196 3596
rect 462280 3556 582196 3584
rect 462280 3544 462286 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 229465 3519 229523 3525
rect 229465 3485 229477 3519
rect 229511 3516 229523 3519
rect 231857 3519 231915 3525
rect 231857 3516 231869 3519
rect 229511 3488 231869 3516
rect 229511 3485 229523 3488
rect 229465 3479 229523 3485
rect 231857 3485 231869 3488
rect 231903 3485 231915 3519
rect 233326 3516 233332 3528
rect 231857 3479 231915 3485
rect 231964 3488 233332 3516
rect 230658 3448 230664 3460
rect 229388 3420 230664 3448
rect 230658 3408 230664 3420
rect 230716 3408 230722 3460
rect 230753 3451 230811 3457
rect 230753 3417 230765 3451
rect 230799 3448 230811 3451
rect 231964 3448 231992 3488
rect 233326 3476 233332 3488
rect 233384 3476 233390 3528
rect 233418 3476 233424 3528
rect 233476 3516 233482 3528
rect 234522 3516 234528 3528
rect 233476 3488 234528 3516
rect 233476 3476 233482 3488
rect 234522 3476 234528 3488
rect 234580 3476 234586 3528
rect 234614 3476 234620 3528
rect 234672 3516 234678 3528
rect 235902 3516 235908 3528
rect 234672 3488 235908 3516
rect 234672 3476 234678 3488
rect 235902 3476 235908 3488
rect 235960 3476 235966 3528
rect 258166 3516 258172 3528
rect 236012 3488 258172 3516
rect 230799 3420 231992 3448
rect 230799 3417 230811 3420
rect 230753 3411 230811 3417
rect 232222 3408 232228 3460
rect 232280 3448 232286 3460
rect 236012 3448 236040 3488
rect 258166 3476 258172 3488
rect 258224 3476 258230 3528
rect 258258 3476 258264 3528
rect 258316 3516 258322 3528
rect 259362 3516 259368 3528
rect 258316 3488 259368 3516
rect 258316 3476 258322 3488
rect 259362 3476 259368 3488
rect 259420 3476 259426 3528
rect 259454 3476 259460 3528
rect 259512 3516 259518 3528
rect 260742 3516 260748 3528
rect 259512 3488 260748 3516
rect 259512 3476 259518 3488
rect 260742 3476 260748 3488
rect 260800 3476 260806 3528
rect 261754 3476 261760 3528
rect 261812 3516 261818 3528
rect 262858 3516 262864 3528
rect 261812 3488 262864 3516
rect 261812 3476 261818 3488
rect 262858 3476 262864 3488
rect 262916 3476 262922 3528
rect 262950 3476 262956 3528
rect 263008 3516 263014 3528
rect 263502 3516 263508 3528
rect 263008 3488 263508 3516
rect 263008 3476 263014 3488
rect 263502 3476 263508 3488
rect 263560 3476 263566 3528
rect 264146 3476 264152 3528
rect 264204 3516 264210 3528
rect 264882 3516 264888 3528
rect 264204 3488 264888 3516
rect 264204 3476 264210 3488
rect 264882 3476 264888 3488
rect 264940 3476 264946 3528
rect 265342 3476 265348 3528
rect 265400 3516 265406 3528
rect 266998 3516 267004 3528
rect 265400 3488 267004 3516
rect 265400 3476 265406 3488
rect 266998 3476 267004 3488
rect 267056 3476 267062 3528
rect 273622 3476 273628 3528
rect 273680 3516 273686 3528
rect 274542 3516 274548 3528
rect 273680 3488 274548 3516
rect 273680 3476 273686 3488
rect 274542 3476 274548 3488
rect 274600 3476 274606 3528
rect 280706 3476 280712 3528
rect 280764 3516 280770 3528
rect 281442 3516 281448 3528
rect 280764 3488 281448 3516
rect 280764 3476 280770 3488
rect 281442 3476 281448 3488
rect 281500 3476 281506 3528
rect 284294 3476 284300 3528
rect 284352 3516 284358 3528
rect 285582 3516 285588 3528
rect 284352 3488 285588 3516
rect 284352 3476 284358 3488
rect 285582 3476 285588 3488
rect 285640 3476 285646 3528
rect 287790 3476 287796 3528
rect 287848 3516 287854 3528
rect 288342 3516 288348 3528
rect 287848 3488 288348 3516
rect 287848 3476 287854 3488
rect 288342 3476 288348 3488
rect 288400 3476 288406 3528
rect 288986 3476 288992 3528
rect 289044 3516 289050 3528
rect 289722 3516 289728 3528
rect 289044 3488 289728 3516
rect 289044 3476 289050 3488
rect 289722 3476 289728 3488
rect 289780 3476 289786 3528
rect 290182 3476 290188 3528
rect 290240 3516 290246 3528
rect 291286 3516 291292 3528
rect 290240 3488 291292 3516
rect 290240 3476 290246 3488
rect 291286 3476 291292 3488
rect 291344 3476 291350 3528
rect 291378 3476 291384 3528
rect 291436 3516 291442 3528
rect 292482 3516 292488 3528
rect 291436 3488 292488 3516
rect 291436 3476 291442 3488
rect 292482 3476 292488 3488
rect 292540 3476 292546 3528
rect 294046 3476 294052 3528
rect 294104 3516 294110 3528
rect 294874 3516 294880 3528
rect 294104 3488 294880 3516
rect 294104 3476 294110 3488
rect 294874 3476 294880 3488
rect 294932 3476 294938 3528
rect 295426 3476 295432 3528
rect 295484 3516 295490 3528
rect 296070 3516 296076 3528
rect 295484 3488 296076 3516
rect 295484 3476 295490 3488
rect 296070 3476 296076 3488
rect 296128 3476 296134 3528
rect 298738 3476 298744 3528
rect 298796 3516 298802 3528
rect 299658 3516 299664 3528
rect 298796 3488 299664 3516
rect 298796 3476 298802 3488
rect 299658 3476 299664 3488
rect 299716 3476 299722 3528
rect 307662 3476 307668 3528
rect 307720 3516 307726 3528
rect 315022 3516 315028 3528
rect 307720 3488 315028 3516
rect 307720 3476 307726 3488
rect 315022 3476 315028 3488
rect 315080 3476 315086 3528
rect 315117 3519 315175 3525
rect 315117 3485 315129 3519
rect 315163 3516 315175 3519
rect 320910 3516 320916 3528
rect 315163 3488 320916 3516
rect 315163 3485 315175 3488
rect 315117 3479 315175 3485
rect 320910 3476 320916 3488
rect 320968 3476 320974 3528
rect 322198 3476 322204 3528
rect 322256 3516 322262 3528
rect 323302 3516 323308 3528
rect 322256 3488 323308 3516
rect 322256 3476 322262 3488
rect 323302 3476 323308 3488
rect 323360 3476 323366 3528
rect 324130 3476 324136 3528
rect 324188 3516 324194 3528
rect 344554 3516 344560 3528
rect 324188 3488 344560 3516
rect 324188 3476 324194 3488
rect 344554 3476 344560 3488
rect 344612 3476 344618 3528
rect 344922 3476 344928 3528
rect 344980 3516 344986 3528
rect 379974 3516 379980 3528
rect 344980 3488 379980 3516
rect 344980 3476 344986 3488
rect 379974 3476 379980 3488
rect 380032 3476 380038 3528
rect 386322 3476 386328 3528
rect 386380 3516 386386 3528
rect 450906 3516 450912 3528
rect 386380 3488 450912 3516
rect 386380 3476 386386 3488
rect 450906 3476 450912 3488
rect 450964 3476 450970 3528
rect 453942 3476 453948 3528
rect 454000 3516 454006 3528
rect 456610 3516 456616 3528
rect 454000 3488 456616 3516
rect 454000 3476 454006 3488
rect 456610 3476 456616 3488
rect 456668 3476 456674 3528
rect 456794 3476 456800 3528
rect 456852 3516 456858 3528
rect 458082 3516 458088 3528
rect 456852 3488 458088 3516
rect 456852 3476 456858 3488
rect 458082 3476 458088 3488
rect 458140 3476 458146 3528
rect 458174 3476 458180 3528
rect 458232 3516 458238 3528
rect 568022 3516 568028 3528
rect 458232 3488 568028 3516
rect 458232 3476 458238 3488
rect 568022 3476 568028 3488
rect 568080 3476 568086 3528
rect 569218 3476 569224 3528
rect 569276 3516 569282 3528
rect 570322 3516 570328 3528
rect 569276 3488 570328 3516
rect 569276 3476 569282 3488
rect 570322 3476 570328 3488
rect 570380 3476 570386 3528
rect 232280 3420 236040 3448
rect 236089 3451 236147 3457
rect 232280 3408 232286 3420
rect 236089 3417 236101 3451
rect 236135 3448 236147 3451
rect 236135 3420 240364 3448
rect 236135 3417 236147 3420
rect 236089 3411 236147 3417
rect 9950 3340 9956 3392
rect 10008 3380 10014 3392
rect 17218 3380 17224 3392
rect 10008 3352 17224 3380
rect 10008 3340 10014 3352
rect 17218 3340 17224 3352
rect 17276 3340 17282 3392
rect 51350 3340 51356 3392
rect 51408 3380 51414 3392
rect 52362 3380 52368 3392
rect 51408 3352 52368 3380
rect 51408 3340 51414 3352
rect 52362 3340 52368 3352
rect 52420 3340 52426 3392
rect 58434 3340 58440 3392
rect 58492 3380 58498 3392
rect 59262 3380 59268 3392
rect 58492 3352 59268 3380
rect 58492 3340 58498 3352
rect 59262 3340 59268 3352
rect 59320 3340 59326 3392
rect 67910 3340 67916 3392
rect 67968 3380 67974 3392
rect 71038 3380 71044 3392
rect 67968 3352 71044 3380
rect 67968 3340 67974 3352
rect 71038 3340 71044 3352
rect 71096 3340 71102 3392
rect 71498 3340 71504 3392
rect 71556 3380 71562 3392
rect 72418 3380 72424 3392
rect 71556 3352 72424 3380
rect 71556 3340 71562 3352
rect 72418 3340 72424 3352
rect 72476 3340 72482 3392
rect 74994 3340 75000 3392
rect 75052 3380 75058 3392
rect 76558 3380 76564 3392
rect 75052 3352 76564 3380
rect 75052 3340 75058 3352
rect 76558 3340 76564 3352
rect 76616 3340 76622 3392
rect 85666 3340 85672 3392
rect 85724 3380 85730 3392
rect 172698 3380 172704 3392
rect 85724 3352 172704 3380
rect 85724 3340 85730 3352
rect 172698 3340 172704 3352
rect 172756 3340 172762 3392
rect 205082 3340 205088 3392
rect 205140 3380 205146 3392
rect 205542 3380 205548 3392
rect 205140 3352 205548 3380
rect 205140 3340 205146 3352
rect 205542 3340 205548 3352
rect 205600 3340 205606 3392
rect 213362 3340 213368 3392
rect 213420 3380 213426 3392
rect 213822 3380 213828 3392
rect 213420 3352 213828 3380
rect 213420 3340 213426 3352
rect 213822 3340 213828 3352
rect 213880 3340 213886 3392
rect 214466 3340 214472 3392
rect 214524 3380 214530 3392
rect 215202 3380 215208 3392
rect 214524 3352 215208 3380
rect 214524 3340 214530 3352
rect 215202 3340 215208 3352
rect 215260 3340 215266 3392
rect 238757 3383 238815 3389
rect 238757 3380 238769 3383
rect 215312 3352 238769 3380
rect 6454 3272 6460 3324
rect 6512 3312 6518 3324
rect 7558 3312 7564 3324
rect 6512 3284 7564 3312
rect 6512 3272 6518 3284
rect 7558 3272 7564 3284
rect 7616 3272 7622 3324
rect 38378 3272 38384 3324
rect 38436 3312 38442 3324
rect 43438 3312 43444 3324
rect 38436 3284 43444 3312
rect 38436 3272 38442 3284
rect 43438 3272 43444 3284
rect 43496 3272 43502 3324
rect 92750 3272 92756 3324
rect 92808 3312 92814 3324
rect 176838 3312 176844 3324
rect 92808 3284 176844 3312
rect 92808 3272 92814 3284
rect 176838 3272 176844 3284
rect 176896 3272 176902 3324
rect 89162 3204 89168 3256
rect 89220 3244 89226 3256
rect 98549 3247 98607 3253
rect 98549 3244 98561 3247
rect 89220 3216 98561 3244
rect 89220 3204 89226 3216
rect 98549 3213 98561 3216
rect 98595 3213 98607 3247
rect 98549 3207 98607 3213
rect 98638 3204 98644 3256
rect 98696 3244 98702 3256
rect 99282 3244 99288 3256
rect 98696 3216 99288 3244
rect 98696 3204 98702 3216
rect 99282 3204 99288 3216
rect 99340 3204 99346 3256
rect 179598 3244 179604 3256
rect 99392 3216 179604 3244
rect 53742 3136 53748 3188
rect 53800 3176 53806 3188
rect 57146 3176 57152 3188
rect 53800 3148 57152 3176
rect 53800 3136 53806 3148
rect 57146 3136 57152 3148
rect 57204 3136 57210 3188
rect 96246 3136 96252 3188
rect 96304 3176 96310 3188
rect 99392 3176 99420 3216
rect 179598 3204 179604 3216
rect 179656 3204 179662 3256
rect 209774 3204 209780 3256
rect 209832 3244 209838 3256
rect 215312 3244 215340 3352
rect 238757 3349 238769 3352
rect 238803 3349 238815 3383
rect 238757 3343 238815 3349
rect 238849 3315 238907 3321
rect 238849 3312 238861 3315
rect 209832 3216 215340 3244
rect 215404 3284 238861 3312
rect 209832 3204 209838 3216
rect 96304 3148 99420 3176
rect 96304 3136 96310 3148
rect 99834 3136 99840 3188
rect 99892 3176 99898 3188
rect 180978 3176 180984 3188
rect 99892 3148 180984 3176
rect 99892 3136 99898 3148
rect 180978 3136 180984 3148
rect 181036 3136 181042 3188
rect 212166 3136 212172 3188
rect 212224 3176 212230 3188
rect 215404 3176 215432 3284
rect 238849 3281 238861 3284
rect 238895 3281 238907 3315
rect 240336 3312 240364 3420
rect 240502 3408 240508 3460
rect 240560 3448 240566 3460
rect 241422 3448 241428 3460
rect 240560 3420 241428 3448
rect 240560 3408 240566 3420
rect 241422 3408 241428 3420
rect 241480 3408 241486 3460
rect 241698 3408 241704 3460
rect 241756 3448 241762 3460
rect 242802 3448 242808 3460
rect 241756 3420 242808 3448
rect 241756 3408 241762 3420
rect 242802 3408 242808 3420
rect 242860 3408 242866 3460
rect 242894 3408 242900 3460
rect 242952 3448 242958 3460
rect 244182 3448 244188 3460
rect 242952 3420 244188 3448
rect 242952 3408 242958 3420
rect 244182 3408 244188 3420
rect 244240 3408 244246 3460
rect 246390 3408 246396 3460
rect 246448 3448 246454 3460
rect 246942 3448 246948 3460
rect 246448 3420 246948 3448
rect 246448 3408 246454 3420
rect 246942 3408 246948 3420
rect 247000 3408 247006 3460
rect 248782 3408 248788 3460
rect 248840 3448 248846 3460
rect 249702 3448 249708 3460
rect 248840 3420 249708 3448
rect 248840 3408 248846 3420
rect 249702 3408 249708 3420
rect 249760 3408 249766 3460
rect 249978 3408 249984 3460
rect 250036 3448 250042 3460
rect 251082 3448 251088 3460
rect 250036 3420 251088 3448
rect 250036 3408 250042 3420
rect 251082 3408 251088 3420
rect 251140 3408 251146 3460
rect 251174 3408 251180 3460
rect 251232 3448 251238 3460
rect 252462 3448 252468 3460
rect 251232 3420 252468 3448
rect 251232 3408 251238 3420
rect 252462 3408 252468 3420
rect 252520 3408 252526 3460
rect 255866 3408 255872 3460
rect 255924 3448 255930 3460
rect 256602 3448 256608 3460
rect 255924 3420 256608 3448
rect 255924 3408 255930 3420
rect 256602 3408 256608 3420
rect 256660 3408 256666 3460
rect 257062 3408 257068 3460
rect 257120 3448 257126 3460
rect 257982 3448 257988 3460
rect 257120 3420 257988 3448
rect 257120 3408 257126 3420
rect 257982 3408 257988 3420
rect 258040 3408 258046 3460
rect 272426 3408 272432 3460
rect 272484 3448 272490 3460
rect 273898 3448 273904 3460
rect 272484 3420 273904 3448
rect 272484 3408 272490 3420
rect 273898 3408 273904 3420
rect 273956 3408 273962 3460
rect 279510 3408 279516 3460
rect 279568 3448 279574 3460
rect 280798 3448 280804 3460
rect 279568 3420 280804 3448
rect 279568 3408 279574 3420
rect 280798 3408 280804 3420
rect 280856 3408 280862 3460
rect 306282 3408 306288 3460
rect 306340 3448 306346 3460
rect 313826 3448 313832 3460
rect 306340 3420 313832 3448
rect 306340 3408 306346 3420
rect 313826 3408 313832 3420
rect 313884 3408 313890 3460
rect 314470 3408 314476 3460
rect 314528 3448 314534 3460
rect 326798 3448 326804 3460
rect 314528 3420 326804 3448
rect 314528 3408 314534 3420
rect 326798 3408 326804 3420
rect 326856 3408 326862 3460
rect 326982 3408 326988 3460
rect 327040 3448 327046 3460
rect 348050 3448 348056 3460
rect 327040 3420 348056 3448
rect 327040 3408 327046 3420
rect 348050 3408 348056 3420
rect 348108 3408 348114 3460
rect 349062 3408 349068 3460
rect 349120 3448 349126 3460
rect 387150 3448 387156 3460
rect 349120 3420 387156 3448
rect 349120 3408 349126 3420
rect 387150 3408 387156 3420
rect 387208 3408 387214 3460
rect 389082 3408 389088 3460
rect 389140 3448 389146 3460
rect 454494 3448 454500 3460
rect 389140 3420 454500 3448
rect 389140 3408 389146 3420
rect 454494 3408 454500 3420
rect 454552 3408 454558 3460
rect 456702 3408 456708 3460
rect 456760 3448 456766 3460
rect 571518 3448 571524 3460
rect 456760 3420 571524 3448
rect 456760 3408 456766 3420
rect 571518 3408 571524 3420
rect 571576 3408 571582 3460
rect 244090 3340 244096 3392
rect 244148 3380 244154 3392
rect 244918 3380 244924 3392
rect 244148 3352 244924 3380
rect 244148 3340 244154 3352
rect 244918 3340 244924 3352
rect 244976 3340 244982 3392
rect 254670 3340 254676 3392
rect 254728 3380 254734 3392
rect 255958 3380 255964 3392
rect 254728 3352 255964 3380
rect 254728 3340 254734 3352
rect 255958 3340 255964 3352
rect 256016 3340 256022 3392
rect 313918 3340 313924 3392
rect 313976 3380 313982 3392
rect 325602 3380 325608 3392
rect 313976 3352 325608 3380
rect 313976 3340 313982 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332502 3340 332508 3392
rect 332560 3380 332566 3392
rect 358722 3380 358728 3392
rect 332560 3352 358728 3380
rect 332560 3340 332566 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 368382 3340 368388 3392
rect 368440 3380 368446 3392
rect 418982 3380 418988 3392
rect 368440 3352 418988 3380
rect 368440 3340 368446 3352
rect 418982 3340 418988 3352
rect 419040 3340 419046 3392
rect 436002 3340 436008 3392
rect 436060 3380 436066 3392
rect 536098 3380 536104 3392
rect 436060 3352 536104 3380
rect 436060 3340 436066 3352
rect 536098 3340 536104 3352
rect 536156 3340 536162 3392
rect 540238 3340 540244 3392
rect 540296 3380 540302 3392
rect 541986 3380 541992 3392
rect 540296 3352 541992 3380
rect 540296 3340 540302 3352
rect 541986 3340 541992 3352
rect 542044 3340 542050 3392
rect 544378 3340 544384 3392
rect 544436 3380 544442 3392
rect 545482 3380 545488 3392
rect 544436 3352 545488 3380
rect 544436 3340 544442 3352
rect 545482 3340 545488 3352
rect 545540 3340 545546 3392
rect 551278 3340 551284 3392
rect 551336 3380 551342 3392
rect 552658 3380 552664 3392
rect 551336 3352 552664 3380
rect 551336 3340 551342 3352
rect 552658 3340 552664 3352
rect 552716 3340 552722 3392
rect 558178 3340 558184 3392
rect 558236 3380 558242 3392
rect 559742 3380 559748 3392
rect 558236 3352 559748 3380
rect 558236 3340 558242 3352
rect 559742 3340 559748 3352
rect 559800 3340 559806 3392
rect 560938 3340 560944 3392
rect 560996 3380 561002 3392
rect 563238 3380 563244 3392
rect 560996 3352 563244 3380
rect 560996 3340 561002 3352
rect 563238 3340 563244 3352
rect 563296 3340 563302 3392
rect 256786 3312 256792 3324
rect 240336 3284 256792 3312
rect 238849 3275 238907 3281
rect 256786 3272 256792 3284
rect 256844 3272 256850 3324
rect 271230 3272 271236 3324
rect 271288 3312 271294 3324
rect 271782 3312 271788 3324
rect 271288 3284 271788 3312
rect 271288 3272 271294 3284
rect 271782 3272 271788 3284
rect 271840 3272 271846 3324
rect 300762 3272 300768 3324
rect 300820 3312 300826 3324
rect 304350 3312 304356 3324
rect 300820 3284 304356 3312
rect 300820 3272 300826 3284
rect 304350 3272 304356 3284
rect 304408 3272 304414 3324
rect 318058 3272 318064 3324
rect 318116 3312 318122 3324
rect 329190 3312 329196 3324
rect 318116 3284 329196 3312
rect 318116 3272 318122 3284
rect 329190 3272 329196 3284
rect 329248 3272 329254 3324
rect 329742 3272 329748 3324
rect 329800 3312 329806 3324
rect 354030 3312 354036 3324
rect 329800 3284 354036 3312
rect 329800 3272 329806 3284
rect 354030 3272 354036 3284
rect 354088 3272 354094 3324
rect 364242 3272 364248 3324
rect 364300 3312 364306 3324
rect 411898 3312 411904 3324
rect 364300 3284 411904 3312
rect 364300 3272 364306 3284
rect 411898 3272 411904 3284
rect 411956 3272 411962 3324
rect 433150 3272 433156 3324
rect 433208 3312 433214 3324
rect 532510 3312 532516 3324
rect 433208 3284 532516 3312
rect 433208 3272 433214 3284
rect 532510 3272 532516 3284
rect 532568 3272 532574 3324
rect 219250 3204 219256 3256
rect 219308 3244 219314 3256
rect 251266 3244 251272 3256
rect 219308 3216 251272 3244
rect 219308 3204 219314 3216
rect 251266 3204 251272 3216
rect 251324 3204 251330 3256
rect 311158 3204 311164 3256
rect 311216 3244 311222 3256
rect 318518 3244 318524 3256
rect 311216 3216 318524 3244
rect 311216 3204 311222 3216
rect 318518 3204 318524 3216
rect 318576 3204 318582 3256
rect 331122 3204 331128 3256
rect 331180 3244 331186 3256
rect 355226 3244 355232 3256
rect 331180 3216 355232 3244
rect 331180 3204 331186 3216
rect 355226 3204 355232 3216
rect 355284 3204 355290 3256
rect 361482 3204 361488 3256
rect 361540 3244 361546 3256
rect 408402 3244 408408 3256
rect 361540 3216 408408 3244
rect 361540 3204 361546 3216
rect 408402 3204 408408 3216
rect 408460 3204 408466 3256
rect 431862 3204 431868 3256
rect 431920 3244 431926 3256
rect 529014 3244 529020 3256
rect 431920 3216 529020 3244
rect 431920 3204 431926 3216
rect 529014 3204 529020 3216
rect 529072 3204 529078 3256
rect 212224 3148 215432 3176
rect 212224 3136 212230 3148
rect 216858 3136 216864 3188
rect 216916 3176 216922 3188
rect 249886 3176 249892 3188
rect 216916 3148 249892 3176
rect 216916 3136 216922 3148
rect 249886 3136 249892 3148
rect 249944 3136 249950 3188
rect 266538 3136 266544 3188
rect 266596 3176 266602 3188
rect 267642 3176 267648 3188
rect 266596 3148 267648 3176
rect 266596 3136 266602 3148
rect 267642 3136 267648 3148
rect 267700 3136 267706 3188
rect 328270 3136 328276 3188
rect 328328 3176 328334 3188
rect 350442 3176 350448 3188
rect 328328 3148 350448 3176
rect 328328 3136 328334 3148
rect 350442 3136 350448 3148
rect 350500 3136 350506 3188
rect 360102 3136 360108 3188
rect 360160 3176 360166 3188
rect 404814 3176 404820 3188
rect 360160 3148 404820 3176
rect 360160 3136 360166 3148
rect 404814 3136 404820 3148
rect 404872 3136 404878 3188
rect 429102 3136 429108 3188
rect 429160 3176 429166 3188
rect 525426 3176 525432 3188
rect 429160 3148 525432 3176
rect 429160 3136 429166 3148
rect 525426 3136 525432 3148
rect 525484 3136 525490 3188
rect 31294 3068 31300 3120
rect 31352 3108 31358 3120
rect 33778 3108 33784 3120
rect 31352 3080 33784 3108
rect 31352 3068 31358 3080
rect 33778 3068 33784 3080
rect 33836 3068 33842 3120
rect 103330 3068 103336 3120
rect 103388 3108 103394 3120
rect 183830 3108 183836 3120
rect 103388 3080 183836 3108
rect 103388 3068 103394 3080
rect 183830 3068 183836 3080
rect 183888 3068 183894 3120
rect 215662 3068 215668 3120
rect 215720 3108 215726 3120
rect 248598 3108 248604 3120
rect 215720 3080 248604 3108
rect 215720 3068 215726 3080
rect 248598 3068 248604 3080
rect 248656 3068 248662 3120
rect 299382 3068 299388 3120
rect 299440 3108 299446 3120
rect 301958 3108 301964 3120
rect 299440 3080 301964 3108
rect 299440 3068 299446 3080
rect 301958 3068 301964 3080
rect 302016 3068 302022 3120
rect 324222 3068 324228 3120
rect 324280 3108 324286 3120
rect 343358 3108 343364 3120
rect 324280 3080 343364 3108
rect 324280 3068 324286 3080
rect 343358 3068 343364 3080
rect 343416 3068 343422 3120
rect 355962 3068 355968 3120
rect 356020 3108 356026 3120
rect 397730 3108 397736 3120
rect 356020 3080 397736 3108
rect 356020 3068 356026 3080
rect 397730 3068 397736 3080
rect 397788 3068 397794 3120
rect 427722 3068 427728 3120
rect 427780 3108 427786 3120
rect 521838 3108 521844 3120
rect 427780 3080 521844 3108
rect 427780 3068 427786 3080
rect 521838 3068 521844 3080
rect 521896 3068 521902 3120
rect 27706 3000 27712 3052
rect 27764 3040 27770 3052
rect 29638 3040 29644 3052
rect 27764 3012 29644 3040
rect 27764 3000 27770 3012
rect 29638 3000 29644 3012
rect 29696 3000 29702 3052
rect 105722 3000 105728 3052
rect 105780 3040 105786 3052
rect 106182 3040 106188 3052
rect 105780 3012 106188 3040
rect 105780 3000 105786 3012
rect 106182 3000 106188 3012
rect 106240 3000 106246 3052
rect 106918 3000 106924 3052
rect 106976 3040 106982 3052
rect 107562 3040 107568 3052
rect 106976 3012 107568 3040
rect 106976 3000 106982 3012
rect 107562 3000 107568 3012
rect 107620 3000 107626 3052
rect 110506 3000 110512 3052
rect 110564 3040 110570 3052
rect 187694 3040 187700 3052
rect 110564 3012 187700 3040
rect 110564 3000 110570 3012
rect 187694 3000 187700 3012
rect 187752 3000 187758 3052
rect 190822 3000 190828 3052
rect 190880 3040 190886 3052
rect 191742 3040 191748 3052
rect 190880 3012 191748 3040
rect 190880 3000 190886 3012
rect 191742 3000 191748 3012
rect 191800 3000 191806 3052
rect 222746 3000 222752 3052
rect 222804 3040 222810 3052
rect 223482 3040 223488 3052
rect 222804 3012 223488 3040
rect 222804 3000 222810 3012
rect 223482 3000 223488 3012
rect 223540 3000 223546 3052
rect 223942 3000 223948 3052
rect 224000 3040 224006 3052
rect 224862 3040 224868 3052
rect 224000 3012 224868 3040
rect 224000 3000 224006 3012
rect 224862 3000 224868 3012
rect 224920 3000 224926 3052
rect 226334 3000 226340 3052
rect 226392 3040 226398 3052
rect 229649 3043 229707 3049
rect 229649 3040 229661 3043
rect 226392 3012 229661 3040
rect 226392 3000 226398 3012
rect 229649 3009 229661 3012
rect 229695 3009 229707 3043
rect 251450 3040 251456 3052
rect 229649 3003 229707 3009
rect 229756 3012 251456 3040
rect 50154 2932 50160 2984
rect 50212 2972 50218 2984
rect 53098 2972 53104 2984
rect 50212 2944 53104 2972
rect 50212 2932 50218 2944
rect 53098 2932 53104 2944
rect 53156 2932 53162 2984
rect 114002 2932 114008 2984
rect 114060 2972 114066 2984
rect 114462 2972 114468 2984
rect 114060 2944 114468 2972
rect 114060 2932 114066 2944
rect 114462 2932 114468 2944
rect 114520 2932 114526 2984
rect 123478 2932 123484 2984
rect 123536 2972 123542 2984
rect 124122 2972 124128 2984
rect 123536 2944 124128 2972
rect 123536 2932 123542 2944
rect 124122 2932 124128 2944
rect 124180 2932 124186 2984
rect 191834 2972 191840 2984
rect 126164 2944 191840 2972
rect 121086 2864 121092 2916
rect 121144 2904 121150 2916
rect 126057 2907 126115 2913
rect 126057 2904 126069 2907
rect 121144 2876 126069 2904
rect 121144 2864 121150 2876
rect 126057 2873 126069 2876
rect 126103 2873 126115 2907
rect 126057 2867 126115 2873
rect 117590 2796 117596 2848
rect 117648 2836 117654 2848
rect 126164 2836 126192 2944
rect 191834 2932 191840 2944
rect 191892 2932 191898 2984
rect 220446 2932 220452 2984
rect 220504 2972 220510 2984
rect 229756 2972 229784 3012
rect 251450 3000 251456 3012
rect 251508 3000 251514 3052
rect 274818 3000 274824 3052
rect 274876 3040 274882 3052
rect 276658 3040 276664 3052
rect 274876 3012 276664 3040
rect 274876 3000 274882 3012
rect 276658 3000 276664 3012
rect 276716 3000 276722 3052
rect 281902 3000 281908 3052
rect 281960 3040 281966 3052
rect 282822 3040 282828 3052
rect 281960 3012 282828 3040
rect 281960 3000 281966 3012
rect 282822 3000 282828 3012
rect 282880 3000 282886 3052
rect 320082 3000 320088 3052
rect 320140 3040 320146 3052
rect 336274 3040 336280 3052
rect 320140 3012 336280 3040
rect 320140 3000 320146 3012
rect 336274 3000 336280 3012
rect 336332 3000 336338 3052
rect 424778 3000 424784 3052
rect 424836 3040 424842 3052
rect 518342 3040 518348 3052
rect 424836 3012 518348 3040
rect 424836 3000 424842 3012
rect 518342 3000 518348 3012
rect 518400 3000 518406 3052
rect 220504 2944 229784 2972
rect 229833 2975 229891 2981
rect 220504 2932 220510 2944
rect 229833 2941 229845 2975
rect 229879 2972 229891 2975
rect 255406 2972 255412 2984
rect 229879 2944 255412 2972
rect 229879 2941 229891 2944
rect 229833 2935 229891 2941
rect 255406 2932 255412 2944
rect 255464 2932 255470 2984
rect 303430 2932 303436 2984
rect 303488 2972 303494 2984
rect 307938 2972 307944 2984
rect 303488 2944 307944 2972
rect 303488 2932 303494 2944
rect 307938 2932 307944 2944
rect 307996 2932 308002 2984
rect 318610 2932 318616 2984
rect 318668 2972 318674 2984
rect 333882 2972 333888 2984
rect 318668 2944 333888 2972
rect 318668 2932 318674 2944
rect 333882 2932 333888 2944
rect 333940 2932 333946 2984
rect 420822 2932 420828 2984
rect 420880 2972 420886 2984
rect 511258 2972 511264 2984
rect 420880 2944 511264 2972
rect 420880 2932 420886 2944
rect 511258 2932 511264 2944
rect 511316 2932 511322 2984
rect 126241 2907 126299 2913
rect 126241 2873 126253 2907
rect 126287 2904 126299 2907
rect 193398 2904 193404 2916
rect 126287 2876 193404 2904
rect 126287 2873 126299 2876
rect 126241 2867 126299 2873
rect 193398 2864 193404 2876
rect 193456 2864 193462 2916
rect 225138 2864 225144 2916
rect 225196 2904 225202 2916
rect 254118 2904 254124 2916
rect 225196 2876 254124 2904
rect 225196 2864 225202 2876
rect 254118 2864 254124 2876
rect 254176 2864 254182 2916
rect 400122 2864 400128 2916
rect 400180 2904 400186 2916
rect 475746 2904 475752 2916
rect 400180 2876 475752 2904
rect 400180 2864 400186 2876
rect 475746 2864 475752 2876
rect 475804 2864 475810 2916
rect 489178 2864 489184 2916
rect 489236 2904 489242 2916
rect 489914 2904 489920 2916
rect 489236 2876 489920 2904
rect 489236 2864 489242 2876
rect 489914 2864 489920 2876
rect 489972 2864 489978 2916
rect 501598 2864 501604 2916
rect 501656 2904 501662 2916
rect 504174 2904 504180 2916
rect 501656 2876 504180 2904
rect 501656 2864 501662 2876
rect 504174 2864 504180 2876
rect 504232 2864 504238 2916
rect 196158 2836 196164 2848
rect 117648 2808 126192 2836
rect 126256 2808 196164 2836
rect 117648 2796 117654 2808
rect 124674 2728 124680 2780
rect 124732 2768 124738 2780
rect 126256 2768 126284 2808
rect 196158 2796 196164 2808
rect 196216 2796 196222 2848
rect 228726 2796 228732 2848
rect 228784 2836 228790 2848
rect 256878 2836 256884 2848
rect 228784 2808 256884 2836
rect 228784 2796 228790 2808
rect 256878 2796 256884 2808
rect 256936 2796 256942 2848
rect 395982 2796 395988 2848
rect 396040 2836 396046 2848
rect 468662 2836 468668 2848
rect 396040 2808 468668 2836
rect 396040 2796 396046 2808
rect 468662 2796 468668 2808
rect 468720 2796 468726 2848
rect 124732 2740 126284 2768
rect 124732 2728 124738 2740
rect 448514 2728 448520 2780
rect 448572 2768 448578 2780
rect 449802 2768 449808 2780
rect 448572 2740 449808 2768
rect 448572 2728 448578 2740
rect 449802 2728 449808 2740
rect 449860 2728 449866 2780
<< via1 >>
rect 154120 700952 154172 701004
rect 317420 700952 317472 701004
rect 137836 700884 137888 700936
rect 314660 700884 314712 700936
rect 271788 700816 271840 700868
rect 462320 700816 462372 700868
rect 274548 700748 274600 700800
rect 478512 700748 478564 700800
rect 89168 700680 89220 700732
rect 327080 700680 327132 700732
rect 72976 700612 73028 700664
rect 324320 700612 324372 700664
rect 262128 700544 262180 700596
rect 527180 700544 527232 700596
rect 264888 700476 264940 700528
rect 543464 700476 543516 700528
rect 40500 700408 40552 700460
rect 329840 700408 329892 700460
rect 24308 700340 24360 700392
rect 335360 700340 335412 700392
rect 8116 700272 8168 700324
rect 332600 700272 332652 700324
rect 282828 700204 282880 700256
rect 413652 700204 413704 700256
rect 280068 700136 280120 700188
rect 397460 700136 397512 700188
rect 202788 700068 202840 700120
rect 306380 700068 306432 700120
rect 218980 700000 219032 700052
rect 309140 700000 309192 700052
rect 292488 699932 292540 699984
rect 348792 699932 348844 699984
rect 289728 699864 289780 699916
rect 332508 699864 332560 699916
rect 267648 699796 267700 699848
rect 296720 699796 296772 699848
rect 283840 699728 283892 699780
rect 299572 699728 299624 699780
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 253848 696940 253900 696992
rect 580172 696940 580224 696992
rect 256608 683204 256660 683256
rect 580172 683204 580224 683256
rect 3424 683136 3476 683188
rect 338120 683136 338172 683188
rect 251088 670760 251140 670812
rect 580172 670760 580224 670812
rect 3516 670692 3568 670744
rect 345020 670692 345072 670744
rect 3424 656888 3476 656940
rect 340880 656888 340932 656940
rect 244188 643084 244240 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 347780 632068 347832 632120
rect 248328 630640 248380 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 353300 618264 353352 618316
rect 241428 616836 241480 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 350540 605820 350592 605872
rect 235816 590656 235868 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 356060 579640 356112 579692
rect 238668 576852 238720 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 362868 565836 362920 565888
rect 232320 563048 232372 563100
rect 579804 563048 579856 563100
rect 247132 561620 247184 561672
rect 248328 561620 248380 561672
rect 250076 561620 250128 561672
rect 251088 561620 251140 561672
rect 253020 561620 253072 561672
rect 253848 561620 253900 561672
rect 270868 561620 270920 561672
rect 271788 561620 271840 561672
rect 273812 561620 273864 561672
rect 274548 561620 274600 561672
rect 288624 561620 288676 561672
rect 289728 561620 289780 561672
rect 291660 561620 291712 561672
rect 292488 561620 292540 561672
rect 294604 561484 294656 561536
rect 299480 561484 299532 561536
rect 235908 561416 235960 561468
rect 303528 561416 303580 561468
rect 285680 561348 285732 561400
rect 364340 561348 364392 561400
rect 171048 561280 171100 561332
rect 312452 561280 312504 561332
rect 276756 561212 276808 561264
rect 429200 561212 429252 561264
rect 106188 561144 106240 561196
rect 321284 561144 321336 561196
rect 267924 561076 267976 561128
rect 494060 561076 494112 561128
rect 211528 561008 211580 561060
rect 486424 561008 486476 561060
rect 259000 560940 259052 560992
rect 558920 560940 558972 560992
rect 202604 560872 202656 560924
rect 485044 560872 485096 560924
rect 193680 560804 193732 560856
rect 483664 560804 483716 560856
rect 184848 560736 184900 560788
rect 482284 560736 482336 560788
rect 175924 560668 175976 560720
rect 479524 560668 479576 560720
rect 167000 560600 167052 560652
rect 475384 560600 475436 560652
rect 29644 560532 29696 560584
rect 398472 560532 398524 560584
rect 32404 560464 32456 560516
rect 407396 560464 407448 560516
rect 33784 560396 33836 560448
rect 416228 560396 416280 560448
rect 35164 560328 35216 560380
rect 425152 560328 425204 560380
rect 36544 560260 36596 560312
rect 434076 560260 434128 560312
rect 205548 559580 205600 559632
rect 468484 559580 468536 559632
rect 115204 559512 115256 559564
rect 380624 559512 380676 559564
rect 196716 559444 196768 559496
rect 467104 559444 467156 559496
rect 122104 559376 122156 559428
rect 395528 559376 395580 559428
rect 190736 559308 190788 559360
rect 497464 559308 497516 559360
rect 108304 559240 108356 559292
rect 422208 559240 422260 559292
rect 172980 559172 173032 559224
rect 490564 559172 490616 559224
rect 155132 559104 155184 559156
rect 472624 559104 472676 559156
rect 83464 559036 83516 559088
rect 428096 559036 428148 559088
rect 169944 558968 169996 559020
rect 522304 558968 522356 559020
rect 4804 558900 4856 558952
rect 410340 558900 410392 558952
rect 214472 558220 214524 558272
rect 462964 558220 463016 558272
rect 187792 558152 187844 558204
rect 465724 558152 465776 558204
rect 178868 558084 178920 558136
rect 464344 558084 464396 558136
rect 123484 558016 123536 558068
rect 412916 558016 412968 558068
rect 199844 557948 199896 558000
rect 500224 557948 500276 558000
rect 79324 557880 79376 557932
rect 386420 557880 386472 557932
rect 119344 557812 119396 557864
rect 430764 557812 430816 557864
rect 182088 557744 182140 557796
rect 493324 557744 493376 557796
rect 164148 557676 164200 557728
rect 489184 557676 489236 557728
rect 128728 557608 128780 557660
rect 471244 557608 471296 557660
rect 11704 557540 11756 557592
rect 418988 557540 419040 557592
rect 359556 557447 359608 557456
rect 161296 557379 161348 557388
rect 161296 557345 161305 557379
rect 161305 557345 161339 557379
rect 161339 557345 161348 557379
rect 161296 557336 161348 557345
rect 208952 557379 209004 557388
rect 208952 557345 208961 557379
rect 208961 557345 208995 557379
rect 208995 557345 209004 557379
rect 208952 557336 209004 557345
rect 217784 557379 217836 557388
rect 217784 557345 217793 557379
rect 217793 557345 217827 557379
rect 217827 557345 217836 557379
rect 217784 557336 217836 557345
rect 3332 557200 3384 557252
rect 220728 557336 220780 557388
rect 223488 557336 223540 557388
rect 359556 557413 359565 557447
rect 359565 557413 359599 557447
rect 359599 557413 359608 557447
rect 359556 557404 359608 557413
rect 365628 557447 365680 557456
rect 365628 557413 365637 557447
rect 365637 557413 365671 557447
rect 365671 557413 365680 557447
rect 365628 557404 365680 557413
rect 368480 557447 368532 557456
rect 368480 557413 368489 557447
rect 368489 557413 368523 557447
rect 368523 557413 368532 557447
rect 368480 557404 368532 557413
rect 371516 557447 371568 557456
rect 371516 557413 371525 557447
rect 371525 557413 371559 557447
rect 371559 557413 371568 557447
rect 371516 557404 371568 557413
rect 374460 557447 374512 557456
rect 374460 557413 374469 557447
rect 374469 557413 374503 557447
rect 374503 557413 374512 557447
rect 374460 557404 374512 557413
rect 377404 557447 377456 557456
rect 377404 557413 377413 557447
rect 377413 557413 377447 557447
rect 377447 557413 377456 557447
rect 377404 557404 377456 557413
rect 383752 557447 383804 557456
rect 383752 557413 383761 557447
rect 383761 557413 383795 557447
rect 383795 557413 383804 557447
rect 383752 557404 383804 557413
rect 389180 557447 389232 557456
rect 389180 557413 389189 557447
rect 389189 557413 389223 557447
rect 389223 557413 389232 557447
rect 389180 557404 389232 557413
rect 392124 557447 392176 557456
rect 392124 557413 392133 557447
rect 392133 557413 392167 557447
rect 392167 557413 392176 557447
rect 392124 557404 392176 557413
rect 401140 557447 401192 557456
rect 401140 557413 401149 557447
rect 401149 557413 401183 557447
rect 401183 557413 401192 557447
rect 401140 557404 401192 557413
rect 404176 557447 404228 557456
rect 404176 557413 404185 557447
rect 404185 557413 404219 557447
rect 404219 557413 404228 557447
rect 404176 557404 404228 557413
rect 226616 557336 226668 557388
rect 229560 557336 229612 557388
rect 580724 557336 580776 557388
rect 580816 557268 580868 557320
rect 580632 557132 580684 557184
rect 580448 557064 580500 557116
rect 3148 556996 3200 557048
rect 580540 556928 580592 556980
rect 4068 556860 4120 556912
rect 3240 556792 3292 556844
rect 3976 556724 4028 556776
rect 580356 556656 580408 556708
rect 3884 556588 3936 556640
rect 3792 556520 3844 556572
rect 3700 556452 3752 556504
rect 3608 556384 3660 556436
rect 3516 556316 3568 556368
rect 3424 556248 3476 556300
rect 580264 556180 580316 556232
rect 2872 463632 2924 463684
rect 115204 463632 115256 463684
rect 462964 458124 463016 458176
rect 580172 458124 580224 458176
rect 486424 419432 486476 419484
rect 580172 419432 580224 419484
rect 468484 405628 468536 405680
rect 579620 405628 579672 405680
rect 3332 398760 3384 398812
rect 79324 398760 79376 398812
rect 500224 379448 500276 379500
rect 580172 379448 580224 379500
rect 485044 365644 485096 365696
rect 580172 365644 580224 365696
rect 3332 358708 3384 358760
rect 29644 358708 29696 358760
rect 467104 353200 467156 353252
rect 580172 353200 580224 353252
rect 3332 346332 3384 346384
rect 122104 346332 122156 346384
rect 497464 325592 497516 325644
rect 579896 325592 579948 325644
rect 483664 313216 483716 313268
rect 580172 313216 580224 313268
rect 3516 306280 3568 306332
rect 32404 306280 32456 306332
rect 465724 299412 465776 299464
rect 579620 299412 579672 299464
rect 493324 273164 493376 273216
rect 579896 273164 579948 273216
rect 2780 267384 2832 267436
rect 4804 267384 4856 267436
rect 482284 259360 482336 259412
rect 579804 259360 579856 259412
rect 3424 255212 3476 255264
rect 33784 255212 33836 255264
rect 464344 245556 464396 245608
rect 580172 245556 580224 245608
rect 3424 241408 3476 241460
rect 123484 241408 123536 241460
rect 490564 233180 490616 233232
rect 580172 233180 580224 233232
rect 479524 219376 479576 219428
rect 579896 219376 579948 219428
rect 3332 215228 3384 215280
rect 11704 215228 11756 215280
rect 522304 206932 522356 206984
rect 580172 206932 580224 206984
rect 3424 202784 3476 202836
rect 35164 202784 35216 202836
rect 489184 193128 489236 193180
rect 580172 193128 580224 193180
rect 3424 188980 3476 189032
rect 108304 188980 108356 189032
rect 475384 179324 475436 179376
rect 579988 179324 580040 179376
rect 3240 164160 3292 164212
rect 83464 164160 83516 164212
rect 472624 153144 472676 153196
rect 580172 153144 580224 153196
rect 3424 150356 3476 150408
rect 36544 150356 36596 150408
rect 107568 148996 107620 149048
rect 186044 148996 186096 149048
rect 191748 148996 191800 149048
rect 234712 148996 234764 149048
rect 241428 148996 241480 149048
rect 263600 148996 263652 149048
rect 270408 148996 270460 149048
rect 280712 148996 280764 149048
rect 372620 148996 372672 149048
rect 374644 148996 374696 149048
rect 406292 148996 406344 149048
rect 485780 148996 485832 149048
rect 104164 148928 104216 148980
rect 183284 148928 183336 148980
rect 187608 148928 187660 148980
rect 232688 148928 232740 148980
rect 235908 148928 235960 148980
rect 260104 148928 260156 148980
rect 260748 148928 260800 148980
rect 274548 148928 274600 148980
rect 347964 148928 348016 148980
rect 385224 148928 385276 148980
rect 410432 148928 410484 148980
rect 492680 148928 492732 148980
rect 93124 148860 93176 148912
rect 177120 148860 177172 148912
rect 177304 148860 177356 148912
rect 181260 148860 181312 148912
rect 184204 148860 184256 148912
rect 229928 148860 229980 148912
rect 238668 148860 238720 148912
rect 262220 148860 262272 148912
rect 264888 148860 264940 148912
rect 276940 148860 276992 148912
rect 277216 148860 277268 148912
rect 284116 148860 284168 148912
rect 349344 148860 349396 148912
rect 388076 148860 388128 148912
rect 420000 148860 420052 148912
rect 504364 148860 504416 148912
rect 75184 148792 75236 148844
rect 166816 148792 166868 148844
rect 173164 148792 173216 148844
rect 223764 148792 223816 148844
rect 237288 148792 237340 148844
rect 261484 148792 261536 148844
rect 262864 148792 262916 148844
rect 275928 148792 275980 148844
rect 351368 148792 351420 148844
rect 389732 148792 389784 148844
rect 413100 148792 413152 148844
rect 497464 148792 497516 148844
rect 35164 148724 35216 148776
rect 135260 148724 135312 148776
rect 154856 148724 154908 148776
rect 157892 148724 157944 148776
rect 166264 148724 166316 148776
rect 218980 148724 219032 148776
rect 234528 148724 234580 148776
rect 259460 148724 259512 148776
rect 263508 148724 263560 148776
rect 276572 148724 276624 148776
rect 276664 148724 276716 148776
rect 283472 148724 283524 148776
rect 352748 148724 352800 148776
rect 393504 148724 393556 148776
rect 414480 148724 414532 148776
rect 499580 148724 499632 148776
rect 22744 148656 22796 148708
rect 124956 148656 125008 148708
rect 155224 148656 155276 148708
rect 213460 148656 213512 148708
rect 231768 148656 231820 148708
rect 258080 148656 258132 148708
rect 259368 148656 259420 148708
rect 273812 148656 273864 148708
rect 274548 148656 274600 148708
rect 282736 148656 282788 148708
rect 356888 148656 356940 148708
rect 400404 148656 400456 148708
rect 409052 148656 409104 148708
rect 410800 148656 410852 148708
rect 417240 148656 417292 148708
rect 502984 148656 503036 148708
rect 25504 148588 25556 148640
rect 131856 148588 131908 148640
rect 144368 148588 144420 148640
rect 203156 148588 203208 148640
rect 227628 148588 227680 148640
rect 256056 148588 256108 148640
rect 260656 148588 260708 148640
rect 275192 148588 275244 148640
rect 277308 148588 277360 148640
rect 284852 148588 284904 148640
rect 370596 148588 370648 148640
rect 414664 148588 414716 148640
rect 418620 148588 418672 148640
rect 506480 148588 506532 148640
rect 14464 148520 14516 148572
rect 124312 148520 124364 148572
rect 147128 148520 147180 148572
rect 207296 148520 207348 148572
rect 223488 148520 223540 148572
rect 253296 148520 253348 148572
rect 253848 148520 253900 148572
rect 271144 148520 271196 148572
rect 271788 148520 271840 148572
rect 281356 148520 281408 148572
rect 328736 148520 328788 148572
rect 352012 148520 352064 148572
rect 356152 148520 356204 148572
rect 357348 148520 357400 148572
rect 360292 148520 360344 148572
rect 406384 148520 406436 148572
rect 422760 148520 422812 148572
rect 514760 148520 514812 148572
rect 18604 148452 18656 148504
rect 133144 148452 133196 148504
rect 133328 148452 133380 148504
rect 199016 148452 199068 148504
rect 224868 148452 224920 148504
rect 253940 148452 253992 148504
rect 256608 148452 256660 148504
rect 272524 148452 272576 148504
rect 273904 148452 273956 148504
rect 282092 148452 282144 148504
rect 322572 148452 322624 148504
rect 338764 148452 338816 148504
rect 347228 148452 347280 148504
rect 377404 148452 377456 148504
rect 378876 148452 378928 148504
rect 425704 148452 425756 148504
rect 428280 148452 428332 148504
rect 522304 148452 522356 148504
rect 11704 148384 11756 148436
rect 128360 148384 128412 148436
rect 133236 148384 133288 148436
rect 200396 148384 200448 148436
rect 213828 148384 213880 148436
rect 247776 148384 247828 148436
rect 249708 148384 249760 148436
rect 268384 148384 268436 148436
rect 268936 148384 268988 148436
rect 279332 148384 279384 148436
rect 286968 148384 287020 148436
rect 290280 148384 290332 148436
rect 326712 148384 326764 148436
rect 349252 148384 349304 148436
rect 364432 148384 364484 148436
rect 413284 148384 413336 148436
rect 430304 148384 430356 148436
rect 526444 148384 526496 148436
rect 7564 148316 7616 148368
rect 127716 148316 127768 148368
rect 129004 148316 129056 148368
rect 198372 148316 198424 148368
rect 205548 148316 205600 148368
rect 242992 148316 243044 148368
rect 244924 148316 244976 148368
rect 265624 148316 265676 148368
rect 267188 148316 267240 148368
rect 277952 148316 278004 148368
rect 311624 148316 311676 148368
rect 322204 148316 322256 148368
rect 330760 148316 330812 148368
rect 356152 148316 356204 148368
rect 368572 148316 368624 148368
rect 418804 148316 418856 148368
rect 432604 148316 432656 148368
rect 432696 148316 432748 148368
rect 530584 148316 530636 148368
rect 111064 148248 111116 148300
rect 187424 148248 187476 148300
rect 195244 148248 195296 148300
rect 236092 148248 236144 148300
rect 242808 148248 242860 148300
rect 264244 148248 264296 148300
rect 269028 148248 269080 148300
rect 280068 148248 280120 148300
rect 402152 148248 402204 148300
rect 478880 148248 478932 148300
rect 114468 148180 114520 148232
rect 190184 148180 190236 148232
rect 196624 148180 196676 148232
rect 225788 148180 225840 148232
rect 228364 148180 228416 148232
rect 240232 148180 240284 148232
rect 246948 148180 247000 148232
rect 267004 148180 267056 148232
rect 267648 148180 267700 148232
rect 278688 148180 278740 148232
rect 398012 148180 398064 148232
rect 471980 148180 472032 148232
rect 119436 148112 119488 148164
rect 191472 148112 191524 148164
rect 198004 148112 198056 148164
rect 236828 148112 236880 148164
rect 244188 148112 244240 148164
rect 264612 148112 264664 148164
rect 402888 148112 402940 148164
rect 475384 148112 475436 148164
rect 115204 148044 115256 148096
rect 116584 147976 116636 148028
rect 155868 147976 155920 148028
rect 122104 147908 122156 147960
rect 151728 147908 151780 147960
rect 170404 148044 170456 148096
rect 221004 148044 221056 148096
rect 240784 148044 240836 148096
rect 250536 148044 250588 148096
rect 252468 148044 252520 148096
rect 269764 148044 269816 148096
rect 393964 148044 394016 148096
rect 465080 148044 465132 148096
rect 162216 147976 162268 148028
rect 210700 147976 210752 148028
rect 251088 147976 251140 148028
rect 268660 147976 268712 148028
rect 278688 147976 278740 148028
rect 285496 147976 285548 148028
rect 387064 147976 387116 148028
rect 390100 147976 390152 148028
rect 401508 147976 401560 148028
rect 468484 147976 468536 148028
rect 170956 147908 171008 147960
rect 255964 147908 256016 147960
rect 271420 147908 271472 147960
rect 280804 147908 280856 147960
rect 286232 147908 286284 147960
rect 389824 147908 389876 147960
rect 456800 147908 456852 147960
rect 150440 147840 150492 147892
rect 153752 147840 153804 147892
rect 257988 147840 258040 147892
rect 273168 147840 273220 147892
rect 281448 147840 281500 147892
rect 286876 147840 286928 147892
rect 377496 147840 377548 147892
rect 436100 147840 436152 147892
rect 208400 147772 208452 147824
rect 209044 147772 209096 147824
rect 219440 147772 219492 147824
rect 220084 147772 220136 147824
rect 253204 147772 253256 147824
rect 266268 147772 266320 147824
rect 282828 147772 282880 147824
rect 287612 147772 287664 147824
rect 200764 147704 200816 147756
rect 204536 147704 204588 147756
rect 250444 147704 250496 147756
rect 262588 147704 262640 147756
rect 285496 147704 285548 147756
rect 289636 147772 289688 147824
rect 301964 147772 302016 147824
rect 306564 147772 306616 147824
rect 308864 147772 308916 147824
rect 311164 147772 311216 147824
rect 337660 147772 337712 147824
rect 342904 147772 342956 147824
rect 385040 147772 385092 147824
rect 429844 147772 429896 147824
rect 434444 147772 434496 147824
rect 467104 147772 467156 147824
rect 288348 147704 288400 147756
rect 291016 147704 291068 147756
rect 297824 147704 297876 147756
rect 298744 147704 298796 147756
rect 301320 147704 301372 147756
rect 305184 147704 305236 147756
rect 309508 147704 309560 147756
rect 310428 147704 310480 147756
rect 313004 147704 313056 147756
rect 313924 147704 313976 147756
rect 315028 147704 315080 147756
rect 318064 147704 318116 147756
rect 332876 147704 332928 147756
rect 334624 147704 334676 147756
rect 337016 147704 337068 147756
rect 340144 147704 340196 147756
rect 343824 147704 343876 147756
rect 345664 147704 345716 147756
rect 389180 147704 389232 147756
rect 123484 147636 123536 147688
rect 125600 147636 125652 147688
rect 106188 147568 106240 147620
rect 185308 147636 185360 147688
rect 191104 147636 191156 147688
rect 193588 147636 193640 147688
rect 202144 147636 202196 147688
rect 203892 147636 203944 147688
rect 209044 147636 209096 147688
rect 211436 147636 211488 147688
rect 220084 147636 220136 147688
rect 221740 147636 221792 147688
rect 224224 147636 224276 147688
rect 225144 147636 225196 147688
rect 232504 147636 232556 147688
rect 234068 147636 234120 147688
rect 285588 147636 285640 147688
rect 288992 147636 289044 147688
rect 289728 147636 289780 147688
rect 291660 147636 291712 147688
rect 297180 147636 297232 147688
rect 298284 147636 298336 147688
rect 298560 147636 298612 147688
rect 299664 147636 299716 147688
rect 299940 147636 299992 147688
rect 302424 147636 302476 147688
rect 302700 147636 302752 147688
rect 303436 147636 303488 147688
rect 305460 147636 305512 147688
rect 306196 147636 306248 147688
rect 306748 147636 306800 147688
rect 307668 147636 307720 147688
rect 308128 147636 308180 147688
rect 309784 147636 309836 147688
rect 310888 147636 310940 147688
rect 311808 147636 311860 147688
rect 312268 147636 312320 147688
rect 313188 147636 313240 147688
rect 313648 147636 313700 147688
rect 314476 147636 314528 147688
rect 316408 147636 316460 147688
rect 317236 147636 317288 147688
rect 317788 147636 317840 147688
rect 318616 147636 318668 147688
rect 319168 147636 319220 147688
rect 320088 147636 320140 147688
rect 320548 147636 320600 147688
rect 321376 147636 321428 147688
rect 321928 147636 321980 147688
rect 322848 147636 322900 147688
rect 323216 147636 323268 147688
rect 324228 147636 324280 147688
rect 324596 147636 324648 147688
rect 325516 147636 325568 147688
rect 325976 147636 326028 147688
rect 326988 147636 327040 147688
rect 327356 147636 327408 147688
rect 328276 147636 328328 147688
rect 330116 147636 330168 147688
rect 331128 147636 331180 147688
rect 331496 147636 331548 147688
rect 332416 147636 332468 147688
rect 334256 147636 334308 147688
rect 335268 147636 335320 147688
rect 335636 147636 335688 147688
rect 336556 147636 336608 147688
rect 338396 147636 338448 147688
rect 339408 147636 339460 147688
rect 339684 147636 339736 147688
rect 340696 147636 340748 147688
rect 341064 147636 341116 147688
rect 342168 147636 342220 147688
rect 342444 147636 342496 147688
rect 343548 147636 343600 147688
rect 345204 147636 345256 147688
rect 346216 147636 346268 147688
rect 346584 147636 346636 147688
rect 347688 147636 347740 147688
rect 350724 147636 350776 147688
rect 351828 147636 351880 147688
rect 352104 147636 352156 147688
rect 353208 147636 353260 147688
rect 353484 147636 353536 147688
rect 354588 147636 354640 147688
rect 354864 147636 354916 147688
rect 355968 147636 356020 147688
rect 357532 147636 357584 147688
rect 358728 147636 358780 147688
rect 358912 147636 358964 147688
rect 360108 147636 360160 147688
rect 361672 147636 361724 147688
rect 362868 147636 362920 147688
rect 363052 147636 363104 147688
rect 364248 147636 364300 147688
rect 365812 147636 365864 147688
rect 367008 147636 367060 147688
rect 367192 147636 367244 147688
rect 368388 147636 368440 147688
rect 369952 147636 370004 147688
rect 371148 147636 371200 147688
rect 371332 147636 371384 147688
rect 372528 147636 372580 147688
rect 374000 147636 374052 147688
rect 375288 147636 375340 147688
rect 375380 147636 375432 147688
rect 376668 147636 376720 147688
rect 376760 147636 376812 147688
rect 378048 147636 378100 147688
rect 378140 147636 378192 147688
rect 379428 147636 379480 147688
rect 379520 147636 379572 147688
rect 380808 147636 380860 147688
rect 380900 147636 380952 147688
rect 382096 147636 382148 147688
rect 382280 147636 382332 147688
rect 383568 147636 383620 147688
rect 383660 147636 383712 147688
rect 384948 147636 385000 147688
rect 386420 147636 386472 147688
rect 387708 147636 387760 147688
rect 387800 147636 387852 147688
rect 389088 147636 389140 147688
rect 391204 147636 391256 147688
rect 392584 147636 392636 147688
rect 396632 147636 396684 147688
rect 397368 147636 397420 147688
rect 400772 147636 400824 147688
rect 401508 147636 401560 147688
rect 403532 147636 403584 147688
rect 404268 147636 404320 147688
rect 404912 147636 404964 147688
rect 411812 147636 411864 147688
rect 412548 147636 412600 147688
rect 415860 147636 415912 147688
rect 416596 147636 416648 147688
rect 421380 147636 421432 147688
rect 422208 147636 422260 147688
rect 424140 147636 424192 147688
rect 426900 147636 426952 147688
rect 427728 147636 427780 147688
rect 429568 147636 429620 147688
rect 430488 147636 430540 147688
rect 430948 147704 431000 147756
rect 431868 147704 431920 147756
rect 433708 147704 433760 147756
rect 434628 147704 434680 147756
rect 435088 147704 435140 147756
rect 436008 147704 436060 147756
rect 437848 147704 437900 147756
rect 438676 147704 438728 147756
rect 439228 147704 439280 147756
rect 440148 147704 440200 147756
rect 441988 147704 442040 147756
rect 442816 147704 442868 147756
rect 443368 147704 443420 147756
rect 444288 147704 444340 147756
rect 446036 147704 446088 147756
rect 447048 147704 447100 147756
rect 447416 147704 447468 147756
rect 448428 147704 448480 147756
rect 450176 147704 450228 147756
rect 451188 147704 451240 147756
rect 451556 147704 451608 147756
rect 452568 147704 452620 147756
rect 454316 147704 454368 147756
rect 455236 147704 455288 147756
rect 455696 147704 455748 147756
rect 456708 147704 456760 147756
rect 458456 147704 458508 147756
rect 459468 147704 459520 147756
rect 459836 147704 459888 147756
rect 460848 147704 460900 147756
rect 464344 147704 464396 147756
rect 461216 147636 461268 147688
rect 462228 147636 462280 147688
rect 483020 147568 483072 147620
rect 99288 147500 99340 147552
rect 177304 147500 177356 147552
rect 410800 147500 410852 147552
rect 490012 147500 490064 147552
rect 95148 147432 95200 147484
rect 178500 147432 178552 147484
rect 416688 147432 416740 147484
rect 501604 147432 501656 147484
rect 88248 147364 88300 147416
rect 175004 147364 175056 147416
rect 426164 147364 426216 147416
rect 520280 147364 520332 147416
rect 59268 147296 59320 147348
rect 154856 147296 154908 147348
rect 436468 147296 436520 147348
rect 538220 147296 538272 147348
rect 62028 147228 62080 147280
rect 159916 147228 159968 147280
rect 438492 147228 438544 147280
rect 540244 147228 540296 147280
rect 52368 147160 52420 147212
rect 150440 147160 150492 147212
rect 440608 147160 440660 147212
rect 544384 147160 544436 147212
rect 43444 147092 43496 147144
rect 146208 147092 146260 147144
rect 442632 147092 442684 147144
rect 547880 147092 547932 147144
rect 47584 147024 47636 147076
rect 150348 147024 150400 147076
rect 362960 147024 363012 147076
rect 409880 147024 409932 147076
rect 444748 147024 444800 147076
rect 551284 147024 551336 147076
rect 29644 146956 29696 147008
rect 140044 146956 140096 147008
rect 367100 146956 367152 147008
rect 416780 146956 416832 147008
rect 454960 146956 455012 147008
rect 569224 146956 569276 147008
rect 21364 146888 21416 146940
rect 134524 146888 134576 146940
rect 374644 146888 374696 146940
rect 427820 146888 427872 146940
rect 457076 146888 457128 146940
rect 572720 146888 572772 146940
rect 113088 146820 113140 146872
rect 188988 146820 189040 146872
rect 179512 146276 179564 146328
rect 180156 146276 180208 146328
rect 183652 146276 183704 146328
rect 184388 146276 184440 146328
rect 196072 146276 196124 146328
rect 196716 146276 196768 146328
rect 201500 146276 201552 146328
rect 202236 146276 202288 146328
rect 216680 146276 216732 146328
rect 217324 146276 217376 146328
rect 222200 146276 222252 146328
rect 222844 146276 222896 146328
rect 226340 146276 226392 146328
rect 226892 146276 226944 146328
rect 124128 146140 124180 146192
rect 195612 146140 195664 146192
rect 76564 146072 76616 146124
rect 167460 146072 167512 146124
rect 65524 146004 65576 146056
rect 157248 146004 157300 146056
rect 71044 145936 71096 145988
rect 163412 145936 163464 145988
rect 393228 145936 393280 145988
rect 463700 145936 463752 145988
rect 50344 145868 50396 145920
rect 148324 145868 148376 145920
rect 404176 145868 404228 145920
rect 481640 145868 481692 145920
rect 53104 145800 53156 145852
rect 153108 145800 153160 145852
rect 448796 145800 448848 145852
rect 558184 145800 558236 145852
rect 39304 145732 39356 145784
rect 144184 145732 144236 145784
rect 446772 145732 446824 145784
rect 556252 145732 556304 145784
rect 32404 145664 32456 145716
rect 137284 145664 137336 145716
rect 244280 145664 244332 145716
rect 244740 145664 244792 145716
rect 450912 145664 450964 145716
rect 560944 145664 560996 145716
rect 33784 145596 33836 145648
rect 142068 145596 142120 145648
rect 452936 145596 452988 145648
rect 565820 145596 565872 145648
rect 17224 145528 17276 145580
rect 129740 145528 129792 145580
rect 390100 145528 390152 145580
rect 452660 145528 452712 145580
rect 459100 145528 459152 145580
rect 574744 145528 574796 145580
rect 168380 144848 168432 144900
rect 169300 144848 169352 144900
rect 72424 144304 72476 144356
rect 165436 144304 165488 144356
rect 68284 144236 68336 144288
rect 161296 144236 161348 144288
rect 57244 144168 57296 144220
rect 155132 144168 155184 144220
rect 408316 144168 408368 144220
rect 489184 144168 489236 144220
rect 138020 142128 138072 142180
rect 138204 142128 138256 142180
rect 140780 142128 140832 142180
rect 140964 142128 141016 142180
rect 245660 142128 245712 142180
rect 245844 142128 245896 142180
rect 256700 142128 256752 142180
rect 256884 142128 256936 142180
rect 119988 141380 120040 141432
rect 191104 141380 191156 141432
rect 3240 137912 3292 137964
rect 119344 137912 119396 137964
rect 3976 91740 4028 91792
rect 123484 91740 123536 91792
rect 397276 33736 397328 33788
rect 470600 33736 470652 33788
rect 471244 33056 471296 33108
rect 580172 33056 580224 33108
rect 345664 25508 345716 25560
rect 378140 25508 378192 25560
rect 161388 18572 161440 18624
rect 216772 18572 216824 18624
rect 340696 18572 340748 18624
rect 371240 18572 371292 18624
rect 412456 18572 412508 18624
rect 496820 18572 496872 18624
rect 180708 17212 180760 17264
rect 227812 17212 227864 17264
rect 383476 17212 383528 17264
rect 445760 17212 445812 17264
rect 137652 15852 137704 15904
rect 202144 15852 202196 15904
rect 215208 15852 215260 15904
rect 248512 15852 248564 15904
rect 339316 15852 339368 15904
rect 370136 15852 370188 15904
rect 395896 15852 395948 15904
rect 467472 15852 467524 15904
rect 177948 14424 178000 14476
rect 226432 14424 226484 14476
rect 429844 14424 429896 14476
rect 448520 14424 448572 14476
rect 413284 13676 413336 13728
rect 414296 13676 414348 13728
rect 151728 13064 151780 13116
rect 209044 13064 209096 13116
rect 415308 13064 415360 13116
rect 501328 13064 501380 13116
rect 133420 11704 133472 11756
rect 200212 11704 200264 11756
rect 375196 11704 375248 11756
rect 432052 11704 432104 11756
rect 54944 10276 54996 10328
rect 116584 10276 116636 10328
rect 169668 10276 169720 10328
rect 220084 10276 220136 10328
rect 419448 10276 419500 10328
rect 508872 10276 508924 10328
rect 156604 9256 156656 9308
rect 214012 9256 214064 9308
rect 153016 9188 153068 9240
rect 212632 9188 212684 9240
rect 142436 9120 142488 9172
rect 205732 9120 205784 9172
rect 145932 9052 145984 9104
rect 208492 9052 208544 9104
rect 95056 8984 95108 9036
rect 178132 8984 178184 9036
rect 60832 8916 60884 8968
rect 158812 8916 158864 8968
rect 161296 8916 161348 8968
rect 216680 8916 216732 8968
rect 343456 8916 343508 8968
rect 377680 8916 377732 8968
rect 378048 8916 378100 8968
rect 435548 8916 435600 8968
rect 116400 8236 116452 8288
rect 119436 8236 119488 8288
rect 174268 8236 174320 8288
rect 224224 8236 224276 8288
rect 169576 8168 169628 8220
rect 222292 8168 222344 8220
rect 158904 8100 158956 8152
rect 215392 8100 215444 8152
rect 147128 8032 147180 8084
rect 208400 8032 208452 8084
rect 138848 7964 138900 8016
rect 200764 7964 200816 8016
rect 425704 7964 425756 8016
rect 439136 7964 439188 8016
rect 140044 7896 140096 7948
rect 204352 7896 204404 7948
rect 414664 7896 414716 7948
rect 424876 7896 424928 7948
rect 432604 7896 432656 7948
rect 456892 7896 456944 7948
rect 468484 7896 468536 7948
rect 478144 7896 478196 7948
rect 135260 7828 135312 7880
rect 201500 7828 201552 7880
rect 382096 7828 382148 7880
rect 442632 7828 442684 7880
rect 464344 7828 464396 7880
rect 517152 7828 517204 7880
rect 134156 7760 134208 7812
rect 201592 7760 201644 7812
rect 392584 7760 392636 7812
rect 460388 7760 460440 7812
rect 467104 7760 467156 7812
rect 534908 7760 534960 7812
rect 130568 7692 130620 7744
rect 198832 7692 198884 7744
rect 400036 7692 400088 7744
rect 474556 7692 474608 7744
rect 80888 7624 80940 7676
rect 115204 7624 115256 7676
rect 126980 7624 127032 7676
rect 197452 7624 197504 7676
rect 334624 7624 334676 7676
rect 359924 7624 359976 7676
rect 407028 7624 407080 7676
rect 487620 7624 487672 7676
rect 47860 7556 47912 7608
rect 122104 7556 122156 7608
rect 125876 7556 125928 7608
rect 196072 7556 196124 7608
rect 196808 7556 196860 7608
rect 237472 7556 237524 7608
rect 358636 7556 358688 7608
rect 403624 7556 403676 7608
rect 411168 7556 411220 7608
rect 494704 7556 494756 7608
rect 129372 6876 129424 6928
rect 133236 6876 133288 6928
rect 124220 6808 124272 6860
rect 580172 6808 580224 6860
rect 97448 6740 97500 6792
rect 179512 6740 179564 6792
rect 398748 6740 398800 6792
rect 473452 6740 473504 6792
rect 84476 6672 84528 6724
rect 172612 6672 172664 6724
rect 404268 6672 404320 6724
rect 481732 6672 481784 6724
rect 77392 6604 77444 6656
rect 168472 6604 168524 6656
rect 405648 6604 405700 6656
rect 485228 6604 485280 6656
rect 70308 6536 70360 6588
rect 164240 6536 164292 6588
rect 342076 6536 342128 6588
rect 375196 6536 375248 6588
rect 408408 6536 408460 6588
rect 488816 6536 488868 6588
rect 66720 6468 66772 6520
rect 161572 6468 161624 6520
rect 346216 6468 346268 6520
rect 381176 6468 381228 6520
rect 409788 6468 409840 6520
rect 492312 6468 492364 6520
rect 63224 6400 63276 6452
rect 160100 6400 160152 6452
rect 183744 6400 183796 6452
rect 230572 6400 230624 6452
rect 346308 6400 346360 6452
rect 382372 6400 382424 6452
rect 412548 6400 412600 6452
rect 495900 6400 495952 6452
rect 59636 6332 59688 6384
rect 157432 6332 157484 6384
rect 179052 6332 179104 6384
rect 227720 6332 227772 6384
rect 350448 6332 350500 6384
rect 389456 6332 389508 6384
rect 413928 6332 413980 6384
rect 499396 6332 499448 6384
rect 56048 6264 56100 6316
rect 155960 6264 156012 6316
rect 177856 6264 177908 6316
rect 226340 6264 226392 6316
rect 353208 6264 353260 6316
rect 393044 6264 393096 6316
rect 416596 6264 416648 6316
rect 502892 6264 502944 6316
rect 52552 6196 52604 6248
rect 153292 6196 153344 6248
rect 173256 6196 173308 6248
rect 223672 6196 223724 6248
rect 357348 6196 357400 6248
rect 400036 6196 400088 6248
rect 418068 6196 418120 6248
rect 506480 6196 506532 6248
rect 48964 6128 49016 6180
rect 151820 6128 151872 6180
rect 170772 6128 170824 6180
rect 222200 6128 222252 6180
rect 354496 6128 354548 6180
rect 396540 6128 396592 6180
rect 422116 6128 422168 6180
rect 513564 6128 513616 6180
rect 101036 6060 101088 6112
rect 182272 6060 182324 6112
rect 401508 6060 401560 6112
rect 476948 6060 477000 6112
rect 104532 5992 104584 6044
rect 183652 5992 183704 6044
rect 397368 5992 397420 6044
rect 469864 5992 469916 6044
rect 108120 5924 108172 5976
rect 186412 5924 186464 5976
rect 394608 5924 394660 5976
rect 466276 5924 466328 5976
rect 111616 5856 111668 5908
rect 187792 5856 187844 5908
rect 393228 5856 393280 5908
rect 462780 5856 462832 5908
rect 115204 5788 115256 5840
rect 190552 5788 190604 5840
rect 118792 5720 118844 5772
rect 191932 5720 191984 5772
rect 122288 5652 122340 5704
rect 194600 5652 194652 5704
rect 504364 5584 504416 5636
rect 510068 5584 510120 5636
rect 91560 5516 91612 5568
rect 93124 5516 93176 5568
rect 102232 5516 102284 5568
rect 104164 5516 104216 5568
rect 109316 5516 109368 5568
rect 111064 5516 111116 5568
rect 406384 5516 406436 5568
rect 407212 5516 407264 5568
rect 475384 5516 475436 5568
rect 480536 5516 480588 5568
rect 497464 5516 497516 5568
rect 498200 5516 498252 5568
rect 502984 5516 503036 5568
rect 505376 5516 505428 5568
rect 44272 5448 44324 5500
rect 149152 5448 149204 5500
rect 189724 5448 189776 5500
rect 232504 5448 232556 5500
rect 371148 5448 371200 5500
rect 423772 5448 423824 5500
rect 435916 5448 435968 5500
rect 537208 5448 537260 5500
rect 40684 5380 40736 5432
rect 146392 5380 146444 5432
rect 186136 5380 186188 5432
rect 231952 5380 232004 5432
rect 372436 5380 372488 5432
rect 427268 5380 427320 5432
rect 440056 5380 440108 5432
rect 544292 5380 544344 5432
rect 37188 5312 37240 5364
rect 145012 5312 145064 5364
rect 166080 5312 166132 5364
rect 219440 5312 219492 5364
rect 375288 5312 375340 5364
rect 430856 5312 430908 5364
rect 442816 5312 442868 5364
rect 547880 5312 547932 5364
rect 33600 5244 33652 5296
rect 142252 5244 142304 5296
rect 164884 5244 164936 5296
rect 219532 5244 219584 5296
rect 376576 5244 376628 5296
rect 434444 5244 434496 5296
rect 444196 5244 444248 5296
rect 551468 5244 551520 5296
rect 30104 5176 30156 5228
rect 140872 5176 140924 5228
rect 149520 5176 149572 5228
rect 162124 5176 162176 5228
rect 162492 5176 162544 5228
rect 218152 5176 218204 5228
rect 379428 5176 379480 5228
rect 437940 5176 437992 5228
rect 447048 5176 447100 5228
rect 554964 5176 555016 5228
rect 26516 5108 26568 5160
rect 139492 5108 139544 5160
rect 157800 5108 157852 5160
rect 215300 5108 215352 5160
rect 325516 5108 325568 5160
rect 345756 5108 345808 5160
rect 380716 5108 380768 5160
rect 441528 5108 441580 5160
rect 448336 5108 448388 5160
rect 558552 5108 558604 5160
rect 21824 5040 21876 5092
rect 136640 5040 136692 5092
rect 151820 5040 151872 5092
rect 211252 5040 211304 5092
rect 342904 5040 342956 5092
rect 368204 5040 368256 5092
rect 383568 5040 383620 5092
rect 445024 5040 445076 5092
rect 451188 5040 451240 5092
rect 562048 5040 562100 5092
rect 17040 4972 17092 5024
rect 12348 4904 12400 4956
rect 131212 4904 131264 4956
rect 8760 4836 8812 4888
rect 128452 4836 128504 4888
rect 4068 4768 4120 4820
rect 125692 4768 125744 4820
rect 155408 4972 155460 5024
rect 213920 4972 213972 5024
rect 218060 4972 218112 5024
rect 240784 4972 240836 5024
rect 340144 4972 340196 5024
rect 367008 4972 367060 5024
rect 387708 4972 387760 5024
rect 452108 4972 452160 5024
rect 452476 4972 452528 5024
rect 565636 4972 565688 5024
rect 148324 4904 148376 4956
rect 209872 4904 209924 4956
rect 221556 4904 221608 4956
rect 252652 4904 252704 4956
rect 336556 4904 336608 4956
rect 364616 4904 364668 4956
rect 384856 4904 384908 4956
rect 448612 4904 448664 4956
rect 455236 4904 455288 4956
rect 569132 4904 569184 4956
rect 131764 4836 131816 4888
rect 133144 4836 133196 4888
rect 136456 4836 136508 4888
rect 144184 4836 144236 4888
rect 144736 4836 144788 4888
rect 207112 4836 207164 4888
rect 210976 4836 211028 4888
rect 245752 4836 245804 4888
rect 335176 4836 335228 4888
rect 363512 4836 363564 4888
rect 377404 4836 377456 4888
rect 384764 4836 384816 4888
rect 388996 4836 389048 4888
rect 133972 4768 134024 4820
rect 141240 4768 141292 4820
rect 205640 4768 205692 4820
rect 207388 4768 207440 4820
rect 244372 4768 244424 4820
rect 321376 4768 321428 4820
rect 338672 4768 338724 4820
rect 342168 4768 342220 4820
rect 374092 4768 374144 4820
rect 390468 4768 390520 4820
rect 459192 4836 459244 4888
rect 459468 4836 459520 4888
rect 576308 4836 576360 4888
rect 455696 4768 455748 4820
rect 456616 4768 456668 4820
rect 572720 4768 572772 4820
rect 65524 4700 65576 4752
rect 161480 4700 161532 4752
rect 175464 4700 175516 4752
rect 196624 4700 196676 4752
rect 203892 4700 203944 4752
rect 241612 4700 241664 4752
rect 368296 4700 368348 4752
rect 420184 4700 420236 4752
rect 438676 4700 438728 4752
rect 540796 4700 540848 4752
rect 73804 4632 73856 4684
rect 75184 4632 75236 4684
rect 72608 4564 72660 4616
rect 165712 4632 165764 4684
rect 200304 4632 200356 4684
rect 228364 4632 228416 4684
rect 364156 4632 364208 4684
rect 413100 4632 413152 4684
rect 431776 4632 431828 4684
rect 69112 4496 69164 4548
rect 162860 4564 162912 4616
rect 366916 4564 366968 4616
rect 416688 4564 416740 4616
rect 434628 4564 434680 4616
rect 76196 4428 76248 4480
rect 167000 4496 167052 4548
rect 360016 4496 360068 4548
rect 406016 4496 406068 4548
rect 427636 4496 427688 4548
rect 523040 4496 523092 4548
rect 533712 4632 533764 4684
rect 530124 4496 530176 4548
rect 79692 4428 79744 4480
rect 169852 4428 169904 4480
rect 362868 4428 362920 4480
rect 409604 4428 409656 4480
rect 430488 4428 430540 4480
rect 526628 4428 526680 4480
rect 83280 4360 83332 4412
rect 171232 4360 171284 4412
rect 355876 4360 355928 4412
rect 398932 4360 398984 4412
rect 426256 4360 426308 4412
rect 519544 4360 519596 4412
rect 86868 4292 86920 4344
rect 173992 4292 174044 4344
rect 358728 4292 358780 4344
rect 402520 4292 402572 4344
rect 423588 4292 423640 4344
rect 515956 4292 516008 4344
rect 90364 4224 90416 4276
rect 175372 4224 175424 4276
rect 194416 4224 194468 4276
rect 198004 4224 198056 4276
rect 354588 4224 354640 4276
rect 395344 4224 395396 4276
rect 422208 4224 422260 4276
rect 512460 4224 512512 4276
rect 7656 4156 7708 4208
rect 11704 4156 11756 4208
rect 128176 4156 128228 4208
rect 129004 4156 129056 4208
rect 143540 4156 143592 4208
rect 146944 4156 146996 4208
rect 154212 4156 154264 4208
rect 155224 4156 155276 4208
rect 163688 4156 163740 4208
rect 166264 4156 166316 4208
rect 167184 4156 167236 4208
rect 170404 4156 170456 4208
rect 171968 4156 172020 4208
rect 173164 4156 173216 4208
rect 182548 4156 182600 4208
rect 184204 4156 184256 4208
rect 193220 4156 193272 4208
rect 195244 4156 195296 4208
rect 338764 4156 338816 4208
rect 342168 4156 342220 4208
rect 389824 4156 389876 4208
rect 391848 4156 391900 4208
rect 418804 4156 418856 4208
rect 421380 4156 421432 4208
rect 522304 4156 522356 4208
rect 524236 4156 524288 4208
rect 526444 4156 526496 4208
rect 527824 4156 527876 4208
rect 530584 4156 530636 4208
rect 531320 4156 531372 4208
rect 15936 4088 15988 4140
rect 18604 4088 18656 4140
rect 45468 4088 45520 4140
rect 47584 4088 47636 4140
rect 93952 4088 94004 4140
rect 95148 4088 95200 4140
rect 175280 4088 175332 4140
rect 208584 4088 208636 4140
rect 244280 4088 244332 4140
rect 296628 4088 296680 4140
rect 297272 4088 297324 4140
rect 303528 4088 303580 4140
rect 309048 4088 309100 4140
rect 315948 4088 316000 4140
rect 330392 4088 330444 4140
rect 332416 4088 332468 4140
rect 357532 4088 357584 4140
rect 365628 4088 365680 4140
rect 415492 4088 415544 4140
rect 424784 4088 424836 4140
rect 424968 4088 425020 4140
rect 437296 4088 437348 4140
rect 539600 4088 539652 4140
rect 574744 4088 574796 4140
rect 577412 4088 577464 4140
rect 64328 4020 64380 4072
rect 68284 4020 68336 4072
rect 82084 4020 82136 4072
rect 171140 4020 171192 4072
rect 206192 4020 206244 4072
rect 242992 4020 243044 4072
rect 317236 4020 317288 4072
rect 331588 4020 331640 4072
rect 333888 4020 333940 4072
rect 361120 4020 361172 4072
rect 372528 4020 372580 4072
rect 426164 4020 426216 4072
rect 440148 4020 440200 4072
rect 543188 4020 543240 4072
rect 41880 3952 41932 4004
rect 50344 3952 50396 4004
rect 57244 3952 57296 4004
rect 65432 3952 65484 4004
rect 78588 3952 78640 4004
rect 168380 3952 168432 4004
rect 201500 3952 201552 4004
rect 46664 3884 46716 3936
rect 150532 3884 150584 3936
rect 202696 3884 202748 3936
rect 241520 3952 241572 4004
rect 307576 3952 307628 4004
rect 318708 3952 318760 4004
rect 247224 3884 247276 3936
rect 310428 3884 310480 3936
rect 319720 3884 319772 3936
rect 332692 3952 332744 4004
rect 335268 3952 335320 4004
rect 362316 3952 362368 4004
rect 369768 3952 369820 4004
rect 422576 3952 422628 4004
rect 441436 3952 441488 4004
rect 546684 3952 546736 4004
rect 335084 3884 335136 3936
rect 336648 3884 336700 3936
rect 365812 3884 365864 3936
rect 373908 3884 373960 3936
rect 429660 3884 429712 3936
rect 444288 3884 444340 3936
rect 550272 3884 550324 3936
rect 34796 3816 34848 3868
rect 39304 3816 39356 3868
rect 43076 3816 43128 3868
rect 147680 3816 147732 3868
rect 199108 3816 199160 3868
rect 229836 3816 229888 3868
rect 231032 3816 231084 3868
rect 231768 3816 231820 3868
rect 237380 3816 237432 3868
rect 240232 3816 240284 3868
rect 309784 3816 309836 3868
rect 317328 3816 317380 3868
rect 317420 3816 317472 3868
rect 319996 3816 320048 3868
rect 337476 3816 337528 3868
rect 339408 3816 339460 3868
rect 369400 3816 369452 3868
rect 376668 3816 376720 3868
rect 433248 3816 433300 3868
rect 445576 3816 445628 3868
rect 553768 3816 553820 3868
rect 23020 3748 23072 3800
rect 32404 3748 32456 3800
rect 35992 3748 36044 3800
rect 143632 3748 143684 3800
rect 197912 3748 197964 3800
rect 238760 3748 238812 3800
rect 245200 3748 245252 3800
rect 253204 3748 253256 3800
rect 283104 3748 283156 3800
rect 287152 3748 287204 3800
rect 304816 3748 304868 3800
rect 310244 3748 310296 3800
rect 311808 3748 311860 3800
rect 322112 3748 322164 3800
rect 322848 3748 322900 3800
rect 340972 3748 341024 3800
rect 343548 3748 343600 3800
rect 376484 3748 376536 3800
rect 380808 3748 380860 3800
rect 440332 3748 440384 3800
rect 448428 3748 448480 3800
rect 557356 3748 557408 3800
rect 19432 3680 19484 3732
rect 35164 3680 35216 3732
rect 39580 3680 39632 3732
rect 146300 3680 146352 3732
rect 192024 3680 192076 3732
rect 32404 3612 32456 3664
rect 142160 3612 142212 3664
rect 195612 3612 195664 3664
rect 226524 3612 226576 3664
rect 572 3544 624 3596
rect 14464 3544 14516 3596
rect 2872 3476 2924 3528
rect 3976 3476 4028 3528
rect 13544 3476 13596 3528
rect 25504 3544 25556 3596
rect 28908 3544 28960 3596
rect 140964 3544 141016 3596
rect 188528 3544 188580 3596
rect 229928 3680 229980 3732
rect 238852 3680 238904 3732
rect 239312 3680 239364 3732
rect 250444 3680 250496 3732
rect 252376 3680 252428 3732
rect 269212 3680 269264 3732
rect 310336 3680 310388 3732
rect 316224 3680 316276 3732
rect 321468 3680 321520 3732
rect 339868 3680 339920 3732
rect 340788 3680 340840 3732
rect 372896 3680 372948 3732
rect 382188 3680 382240 3732
rect 443828 3680 443880 3732
rect 449716 3680 449768 3732
rect 560852 3680 560904 3732
rect 229836 3612 229888 3664
rect 238116 3612 238168 3664
rect 238668 3612 238720 3664
rect 245844 3612 245896 3664
rect 247592 3612 247644 3664
rect 266452 3612 266504 3664
rect 304908 3612 304960 3664
rect 311440 3612 311492 3664
rect 313188 3612 313240 3664
rect 324412 3612 324464 3664
rect 325608 3612 325660 3664
rect 346952 3612 347004 3664
rect 347688 3612 347740 3664
rect 383568 3612 383620 3664
rect 384948 3612 385000 3664
rect 447416 3612 447468 3664
rect 452568 3612 452620 3664
rect 564440 3612 564492 3664
rect 18236 3476 18288 3528
rect 21364 3476 21416 3528
rect 25320 3476 25372 3528
rect 138112 3476 138164 3528
rect 150624 3476 150676 3528
rect 151728 3476 151780 3528
rect 160100 3476 160152 3528
rect 161388 3476 161440 3528
rect 168380 3476 168432 3528
rect 169668 3476 169720 3528
rect 176660 3476 176712 3528
rect 177948 3476 178000 3528
rect 180248 3476 180300 3528
rect 180708 3476 180760 3528
rect 184940 3476 184992 3528
rect 226524 3476 226576 3528
rect 1676 3408 1728 3460
rect 22744 3408 22796 3460
rect 24216 3408 24268 3460
rect 138204 3408 138256 3460
rect 181444 3408 181496 3460
rect 229284 3408 229336 3460
rect 234712 3544 234764 3596
rect 235816 3544 235868 3596
rect 260932 3544 260984 3596
rect 267740 3544 267792 3596
rect 268936 3544 268988 3596
rect 276020 3544 276072 3596
rect 277216 3544 277268 3596
rect 306196 3544 306248 3596
rect 312636 3544 312688 3596
rect 314568 3544 314620 3596
rect 328000 3544 328052 3596
rect 328368 3544 328420 3596
rect 351644 3544 351696 3596
rect 351828 3544 351880 3596
rect 390652 3544 390704 3596
rect 391756 3544 391808 3596
rect 461584 3544 461636 3596
rect 462228 3544 462280 3596
rect 582196 3544 582248 3596
rect 230664 3408 230716 3460
rect 233332 3476 233384 3528
rect 233424 3476 233476 3528
rect 234528 3476 234580 3528
rect 234620 3476 234672 3528
rect 235908 3476 235960 3528
rect 232228 3408 232280 3460
rect 258172 3476 258224 3528
rect 258264 3476 258316 3528
rect 259368 3476 259420 3528
rect 259460 3476 259512 3528
rect 260748 3476 260800 3528
rect 261760 3476 261812 3528
rect 262864 3476 262916 3528
rect 262956 3476 263008 3528
rect 263508 3476 263560 3528
rect 264152 3476 264204 3528
rect 264888 3476 264940 3528
rect 265348 3476 265400 3528
rect 267004 3476 267056 3528
rect 273628 3476 273680 3528
rect 274548 3476 274600 3528
rect 280712 3476 280764 3528
rect 281448 3476 281500 3528
rect 284300 3476 284352 3528
rect 285588 3476 285640 3528
rect 287796 3476 287848 3528
rect 288348 3476 288400 3528
rect 288992 3476 289044 3528
rect 289728 3476 289780 3528
rect 290188 3476 290240 3528
rect 291292 3476 291344 3528
rect 291384 3476 291436 3528
rect 292488 3476 292540 3528
rect 294052 3476 294104 3528
rect 294880 3476 294932 3528
rect 295432 3476 295484 3528
rect 296076 3476 296128 3528
rect 298744 3476 298796 3528
rect 299664 3476 299716 3528
rect 307668 3476 307720 3528
rect 315028 3476 315080 3528
rect 320916 3476 320968 3528
rect 322204 3476 322256 3528
rect 323308 3476 323360 3528
rect 324136 3476 324188 3528
rect 344560 3476 344612 3528
rect 344928 3476 344980 3528
rect 379980 3476 380032 3528
rect 386328 3476 386380 3528
rect 450912 3476 450964 3528
rect 453948 3476 454000 3528
rect 456616 3476 456668 3528
rect 456800 3476 456852 3528
rect 458088 3476 458140 3528
rect 458180 3476 458232 3528
rect 568028 3476 568080 3528
rect 569224 3476 569276 3528
rect 570328 3476 570380 3528
rect 9956 3340 10008 3392
rect 17224 3340 17276 3392
rect 51356 3340 51408 3392
rect 52368 3340 52420 3392
rect 58440 3340 58492 3392
rect 59268 3340 59320 3392
rect 67916 3340 67968 3392
rect 71044 3340 71096 3392
rect 71504 3340 71556 3392
rect 72424 3340 72476 3392
rect 75000 3340 75052 3392
rect 76564 3340 76616 3392
rect 85672 3340 85724 3392
rect 172704 3340 172756 3392
rect 205088 3340 205140 3392
rect 205548 3340 205600 3392
rect 213368 3340 213420 3392
rect 213828 3340 213880 3392
rect 214472 3340 214524 3392
rect 215208 3340 215260 3392
rect 6460 3272 6512 3324
rect 7564 3272 7616 3324
rect 38384 3272 38436 3324
rect 43444 3272 43496 3324
rect 92756 3272 92808 3324
rect 176844 3272 176896 3324
rect 89168 3204 89220 3256
rect 98644 3204 98696 3256
rect 99288 3204 99340 3256
rect 53748 3136 53800 3188
rect 57152 3136 57204 3188
rect 96252 3136 96304 3188
rect 179604 3204 179656 3256
rect 209780 3204 209832 3256
rect 99840 3136 99892 3188
rect 180984 3136 181036 3188
rect 212172 3136 212224 3188
rect 240508 3408 240560 3460
rect 241428 3408 241480 3460
rect 241704 3408 241756 3460
rect 242808 3408 242860 3460
rect 242900 3408 242952 3460
rect 244188 3408 244240 3460
rect 246396 3408 246448 3460
rect 246948 3408 247000 3460
rect 248788 3408 248840 3460
rect 249708 3408 249760 3460
rect 249984 3408 250036 3460
rect 251088 3408 251140 3460
rect 251180 3408 251232 3460
rect 252468 3408 252520 3460
rect 255872 3408 255924 3460
rect 256608 3408 256660 3460
rect 257068 3408 257120 3460
rect 257988 3408 258040 3460
rect 272432 3408 272484 3460
rect 273904 3408 273956 3460
rect 279516 3408 279568 3460
rect 280804 3408 280856 3460
rect 306288 3408 306340 3460
rect 313832 3408 313884 3460
rect 314476 3408 314528 3460
rect 326804 3408 326856 3460
rect 326988 3408 327040 3460
rect 348056 3408 348108 3460
rect 349068 3408 349120 3460
rect 387156 3408 387208 3460
rect 389088 3408 389140 3460
rect 454500 3408 454552 3460
rect 456708 3408 456760 3460
rect 571524 3408 571576 3460
rect 244096 3340 244148 3392
rect 244924 3340 244976 3392
rect 254676 3340 254728 3392
rect 255964 3340 256016 3392
rect 313924 3340 313976 3392
rect 325608 3340 325660 3392
rect 332508 3340 332560 3392
rect 358728 3340 358780 3392
rect 368388 3340 368440 3392
rect 418988 3340 419040 3392
rect 436008 3340 436060 3392
rect 536104 3340 536156 3392
rect 540244 3340 540296 3392
rect 541992 3340 542044 3392
rect 544384 3340 544436 3392
rect 545488 3340 545540 3392
rect 551284 3340 551336 3392
rect 552664 3340 552716 3392
rect 558184 3340 558236 3392
rect 559748 3340 559800 3392
rect 560944 3340 560996 3392
rect 563244 3340 563296 3392
rect 256792 3272 256844 3324
rect 271236 3272 271288 3324
rect 271788 3272 271840 3324
rect 300768 3272 300820 3324
rect 304356 3272 304408 3324
rect 318064 3272 318116 3324
rect 329196 3272 329248 3324
rect 329748 3272 329800 3324
rect 354036 3272 354088 3324
rect 364248 3272 364300 3324
rect 411904 3272 411956 3324
rect 433156 3272 433208 3324
rect 532516 3272 532568 3324
rect 219256 3204 219308 3256
rect 251272 3204 251324 3256
rect 311164 3204 311216 3256
rect 318524 3204 318576 3256
rect 331128 3204 331180 3256
rect 355232 3204 355284 3256
rect 361488 3204 361540 3256
rect 408408 3204 408460 3256
rect 431868 3204 431920 3256
rect 529020 3204 529072 3256
rect 216864 3136 216916 3188
rect 249892 3136 249944 3188
rect 266544 3136 266596 3188
rect 267648 3136 267700 3188
rect 328276 3136 328328 3188
rect 350448 3136 350500 3188
rect 360108 3136 360160 3188
rect 404820 3136 404872 3188
rect 429108 3136 429160 3188
rect 525432 3136 525484 3188
rect 31300 3068 31352 3120
rect 33784 3068 33836 3120
rect 103336 3068 103388 3120
rect 183836 3068 183888 3120
rect 215668 3068 215720 3120
rect 248604 3068 248656 3120
rect 299388 3068 299440 3120
rect 301964 3068 302016 3120
rect 324228 3068 324280 3120
rect 343364 3068 343416 3120
rect 355968 3068 356020 3120
rect 397736 3068 397788 3120
rect 427728 3068 427780 3120
rect 521844 3068 521896 3120
rect 27712 3000 27764 3052
rect 29644 3000 29696 3052
rect 105728 3000 105780 3052
rect 106188 3000 106240 3052
rect 106924 3000 106976 3052
rect 107568 3000 107620 3052
rect 110512 3000 110564 3052
rect 187700 3000 187752 3052
rect 190828 3000 190880 3052
rect 191748 3000 191800 3052
rect 222752 3000 222804 3052
rect 223488 3000 223540 3052
rect 223948 3000 224000 3052
rect 224868 3000 224920 3052
rect 226340 3000 226392 3052
rect 50160 2932 50212 2984
rect 53104 2932 53156 2984
rect 114008 2932 114060 2984
rect 114468 2932 114520 2984
rect 123484 2932 123536 2984
rect 124128 2932 124180 2984
rect 121092 2864 121144 2916
rect 117596 2796 117648 2848
rect 191840 2932 191892 2984
rect 220452 2932 220504 2984
rect 251456 3000 251508 3052
rect 274824 3000 274876 3052
rect 276664 3000 276716 3052
rect 281908 3000 281960 3052
rect 282828 3000 282880 3052
rect 320088 3000 320140 3052
rect 336280 3000 336332 3052
rect 424784 3000 424836 3052
rect 518348 3000 518400 3052
rect 255412 2932 255464 2984
rect 303436 2932 303488 2984
rect 307944 2932 307996 2984
rect 318616 2932 318668 2984
rect 333888 2932 333940 2984
rect 420828 2932 420880 2984
rect 511264 2932 511316 2984
rect 193404 2864 193456 2916
rect 225144 2864 225196 2916
rect 254124 2864 254176 2916
rect 400128 2864 400180 2916
rect 475752 2864 475804 2916
rect 489184 2864 489236 2916
rect 489920 2864 489972 2916
rect 501604 2864 501656 2916
rect 504180 2864 504232 2916
rect 124680 2728 124732 2780
rect 196164 2796 196216 2848
rect 228732 2796 228784 2848
rect 256884 2796 256936 2848
rect 395988 2796 396040 2848
rect 468668 2796 468720 2848
rect 448520 2728 448572 2780
rect 449808 2728 449860 2780
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 40512 700466 40540 703520
rect 72988 700670 73016 703520
rect 89180 700738 89208 703520
rect 89168 700732 89220 700738
rect 89168 700674 89220 700680
rect 72976 700664 73028 700670
rect 72976 700606 73028 700612
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 105464 699718 105492 703520
rect 137848 700942 137876 703520
rect 154132 701010 154160 703520
rect 154120 701004 154172 701010
rect 154120 700946 154172 700952
rect 137836 700936 137888 700942
rect 137836 700878 137888 700884
rect 170324 699718 170352 703520
rect 202800 700126 202828 703520
rect 202788 700120 202840 700126
rect 202788 700062 202840 700068
rect 218992 700058 219020 703520
rect 218980 700052 219032 700058
rect 218980 699994 219032 700000
rect 235184 699718 235212 703520
rect 262128 700596 262180 700602
rect 262128 700538 262180 700544
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 106200 561202 106228 699654
rect 171060 561338 171088 699654
rect 235816 590708 235868 590714
rect 235816 590650 235868 590656
rect 235828 567194 235856 590650
rect 235736 567166 235856 567194
rect 232320 563100 232372 563106
rect 232320 563042 232372 563048
rect 171048 561332 171100 561338
rect 171048 561274 171100 561280
rect 106188 561196 106240 561202
rect 106188 561138 106240 561144
rect 211528 561060 211580 561066
rect 211528 561002 211580 561008
rect 202604 560924 202656 560930
rect 202604 560866 202656 560872
rect 193680 560856 193732 560862
rect 193680 560798 193732 560804
rect 184848 560788 184900 560794
rect 184848 560730 184900 560736
rect 175924 560720 175976 560726
rect 175924 560662 175976 560668
rect 167000 560652 167052 560658
rect 167000 560594 167052 560600
rect 29644 560584 29696 560590
rect 29644 560526 29696 560532
rect 4804 558952 4856 558958
rect 4804 558894 4856 558900
rect 3332 557252 3384 557258
rect 3332 557194 3384 557200
rect 3148 557048 3200 557054
rect 3148 556990 3200 556996
rect 3160 547874 3188 556990
rect 3240 556844 3292 556850
rect 3240 556786 3292 556792
rect 3252 552378 3280 556786
rect 3344 553897 3372 557194
rect 4068 556912 4120 556918
rect 4068 556854 4120 556860
rect 3976 556776 4028 556782
rect 3976 556718 4028 556724
rect 3884 556640 3936 556646
rect 3884 556582 3936 556588
rect 3792 556572 3844 556578
rect 3792 556514 3844 556520
rect 3700 556504 3752 556510
rect 3700 556446 3752 556452
rect 3608 556436 3660 556442
rect 3608 556378 3660 556384
rect 3516 556368 3568 556374
rect 3516 556310 3568 556316
rect 3424 556300 3476 556306
rect 3424 556242 3476 556248
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3252 552350 3372 552378
rect 3160 547846 3280 547874
rect 3252 527921 3280 547846
rect 3238 527912 3294 527921
rect 3238 527847 3294 527856
rect 3344 514865 3372 552350
rect 3330 514856 3386 514865
rect 3330 514791 3386 514800
rect 2872 463684 2924 463690
rect 2872 463626 2924 463632
rect 2884 462641 2912 463626
rect 2870 462632 2926 462641
rect 2870 462567 2926 462576
rect 3332 398812 3384 398818
rect 3332 398754 3384 398760
rect 3344 397497 3372 398754
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3332 346384 3384 346390
rect 3332 346326 3384 346332
rect 3344 345409 3372 346326
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3436 293185 3464 556242
rect 3528 319297 3556 556310
rect 3620 371385 3648 556378
rect 3712 410553 3740 556446
rect 3804 423609 3832 556514
rect 3896 449585 3924 556582
rect 3988 475697 4016 556718
rect 4080 501809 4108 556854
rect 4066 501800 4122 501809
rect 4066 501735 4122 501744
rect 3974 475688 4030 475697
rect 3974 475623 4030 475632
rect 3882 449576 3938 449585
rect 3882 449511 3938 449520
rect 3790 423600 3846 423609
rect 3790 423535 3846 423544
rect 3698 410544 3754 410553
rect 3698 410479 3754 410488
rect 3606 371376 3662 371385
rect 3606 371311 3662 371320
rect 3514 319288 3570 319297
rect 3514 319223 3570 319232
rect 3516 306332 3568 306338
rect 3516 306274 3568 306280
rect 3528 306241 3556 306274
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 4816 267442 4844 558894
rect 11704 557592 11756 557598
rect 11704 557534 11756 557540
rect 2780 267436 2832 267442
rect 2780 267378 2832 267384
rect 4804 267436 4856 267442
rect 4804 267378 4856 267384
rect 2792 267209 2820 267378
rect 2778 267200 2834 267209
rect 2778 267135 2834 267144
rect 3424 255264 3476 255270
rect 3424 255206 3476 255212
rect 3436 254153 3464 255206
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3424 241460 3476 241466
rect 3424 241402 3476 241408
rect 3436 241097 3464 241402
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 11716 215286 11744 557534
rect 29656 358766 29684 560526
rect 32404 560516 32456 560522
rect 32404 560458 32456 560464
rect 29644 358760 29696 358766
rect 29644 358702 29696 358708
rect 32416 306338 32444 560458
rect 33784 560448 33836 560454
rect 33784 560390 33836 560396
rect 32404 306332 32456 306338
rect 32404 306274 32456 306280
rect 33796 255270 33824 560390
rect 35164 560380 35216 560386
rect 35164 560322 35216 560328
rect 33784 255264 33836 255270
rect 33784 255206 33836 255212
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 11704 215280 11756 215286
rect 11704 215222 11756 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 35176 202842 35204 560322
rect 36544 560312 36596 560318
rect 36544 560254 36596 560260
rect 3424 202836 3476 202842
rect 3424 202778 3476 202784
rect 35164 202836 35216 202842
rect 35164 202778 35216 202784
rect 3436 201929 3464 202778
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 36556 150414 36584 560254
rect 115204 559564 115256 559570
rect 115204 559506 115256 559512
rect 108304 559292 108356 559298
rect 108304 559234 108356 559240
rect 83464 559088 83516 559094
rect 83464 559030 83516 559036
rect 79324 557932 79376 557938
rect 79324 557874 79376 557880
rect 79336 398818 79364 557874
rect 79324 398812 79376 398818
rect 79324 398754 79376 398760
rect 83476 164218 83504 559030
rect 108316 189038 108344 559234
rect 115216 463690 115244 559506
rect 122104 559428 122156 559434
rect 122104 559370 122156 559376
rect 119344 557864 119396 557870
rect 119344 557806 119396 557812
rect 115204 463684 115256 463690
rect 115204 463626 115256 463632
rect 108304 189032 108356 189038
rect 108304 188974 108356 188980
rect 83464 164212 83516 164218
rect 83464 164154 83516 164160
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 36544 150408 36596 150414
rect 36544 150350 36596 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 107568 149048 107620 149054
rect 107568 148990 107620 148996
rect 104164 148980 104216 148986
rect 104164 148922 104216 148928
rect 93124 148912 93176 148918
rect 93124 148854 93176 148860
rect 75184 148844 75236 148850
rect 75184 148786 75236 148792
rect 35164 148776 35216 148782
rect 35164 148718 35216 148724
rect 22744 148708 22796 148714
rect 22744 148650 22796 148656
rect 14464 148572 14516 148578
rect 14464 148514 14516 148520
rect 11704 148436 11756 148442
rect 11704 148378 11756 148384
rect 7564 148368 7616 148374
rect 7564 148310 7616 148316
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3422 111752 3478 111761
rect 3422 111687 3478 111696
rect 3436 110673 3464 111687
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3976 91792 4028 91798
rect 3976 91734 4028 91740
rect 3422 85504 3478 85513
rect 3422 85439 3478 85448
rect 3436 84697 3464 85439
rect 3422 84688 3478 84697
rect 3422 84623 3478 84632
rect 3330 59256 3386 59265
rect 3330 59191 3386 59200
rect 3344 58585 3372 59191
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 3330 33144 3386 33153
rect 3330 33079 3386 33088
rect 3344 32473 3372 33079
rect 3330 32464 3386 32473
rect 3330 32399 3386 32408
rect 3422 20632 3478 20641
rect 3422 20567 3478 20576
rect 3436 19417 3464 20567
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 572 3596 624 3602
rect 572 3538 624 3544
rect 584 480 612 3538
rect 3988 3534 4016 91734
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 480 1716 3402
rect 2884 480 2912 3470
rect 4080 480 4108 4762
rect 5262 3360 5318 3369
rect 7576 3330 7604 148310
rect 8760 4888 8812 4894
rect 8760 4830 8812 4836
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 5262 3295 5318 3304
rect 6460 3324 6512 3330
rect 5276 480 5304 3295
rect 6460 3266 6512 3272
rect 7564 3324 7616 3330
rect 7564 3266 7616 3272
rect 6472 480 6500 3266
rect 7668 480 7696 4150
rect 8772 480 8800 4830
rect 11716 4214 11744 148378
rect 12348 4956 12400 4962
rect 12348 4898 12400 4904
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 11150 3496 11206 3505
rect 11150 3431 11206 3440
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9968 480 9996 3334
rect 11164 480 11192 3431
rect 12360 480 12388 4898
rect 14476 3602 14504 148514
rect 18604 148504 18656 148510
rect 18604 148446 18656 148452
rect 17224 145580 17276 145586
rect 17224 145522 17276 145528
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 14738 3632 14794 3641
rect 14464 3596 14516 3602
rect 14738 3567 14794 3576
rect 14464 3538 14516 3544
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13556 480 13584 3470
rect 14752 480 14780 3567
rect 15948 480 15976 4082
rect 17052 480 17080 4966
rect 17236 3398 17264 145522
rect 18616 4146 18644 148446
rect 21364 146940 21416 146946
rect 21364 146882 21416 146888
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 20626 3768 20682 3777
rect 19432 3732 19484 3738
rect 20626 3703 20682 3712
rect 19432 3674 19484 3680
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 18248 480 18276 3470
rect 19444 480 19472 3674
rect 20640 480 20668 3703
rect 21376 3534 21404 146882
rect 21824 5092 21876 5098
rect 21824 5034 21876 5040
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21836 480 21864 5034
rect 22756 3466 22784 148650
rect 25504 148640 25556 148646
rect 25504 148582 25556 148588
rect 23020 3800 23072 3806
rect 23020 3742 23072 3748
rect 22744 3460 22796 3466
rect 22744 3402 22796 3408
rect 23032 480 23060 3742
rect 25516 3602 25544 148582
rect 29644 147008 29696 147014
rect 29644 146950 29696 146956
rect 26516 5160 26568 5166
rect 26516 5102 26568 5108
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 480 24256 3402
rect 25332 480 25360 3470
rect 26528 480 26556 5102
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 27724 480 27752 2994
rect 28920 480 28948 3538
rect 29656 3058 29684 146950
rect 32404 145716 32456 145722
rect 32404 145658 32456 145664
rect 30104 5228 30156 5234
rect 30104 5170 30156 5176
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 30116 480 30144 5170
rect 32416 3806 32444 145658
rect 33784 145648 33836 145654
rect 33784 145590 33836 145596
rect 33600 5296 33652 5302
rect 33600 5238 33652 5244
rect 32404 3800 32456 3806
rect 32404 3742 32456 3748
rect 32404 3664 32456 3670
rect 32404 3606 32456 3612
rect 31300 3120 31352 3126
rect 31300 3062 31352 3068
rect 31312 480 31340 3062
rect 32416 480 32444 3606
rect 33612 480 33640 5238
rect 33796 3126 33824 145590
rect 34796 3868 34848 3874
rect 34796 3810 34848 3816
rect 33784 3120 33836 3126
rect 33784 3062 33836 3068
rect 34808 480 34836 3810
rect 35176 3738 35204 148718
rect 59268 147348 59320 147354
rect 59268 147290 59320 147296
rect 52368 147212 52420 147218
rect 52368 147154 52420 147160
rect 43444 147144 43496 147150
rect 43444 147086 43496 147092
rect 39304 145784 39356 145790
rect 39304 145726 39356 145732
rect 37188 5364 37240 5370
rect 37188 5306 37240 5312
rect 35992 3800 36044 3806
rect 35992 3742 36044 3748
rect 35164 3732 35216 3738
rect 35164 3674 35216 3680
rect 36004 480 36032 3742
rect 37200 480 37228 5306
rect 39316 3874 39344 145726
rect 40684 5432 40736 5438
rect 40684 5374 40736 5380
rect 39304 3868 39356 3874
rect 39304 3810 39356 3816
rect 39580 3732 39632 3738
rect 39580 3674 39632 3680
rect 38384 3324 38436 3330
rect 38384 3266 38436 3272
rect 38396 480 38424 3266
rect 39592 480 39620 3674
rect 40696 480 40724 5374
rect 41880 4004 41932 4010
rect 41880 3946 41932 3952
rect 41892 480 41920 3946
rect 43076 3868 43128 3874
rect 43076 3810 43128 3816
rect 43088 480 43116 3810
rect 43456 3330 43484 147086
rect 47584 147076 47636 147082
rect 47584 147018 47636 147024
rect 44272 5500 44324 5506
rect 44272 5442 44324 5448
rect 43444 3324 43496 3330
rect 43444 3266 43496 3272
rect 44284 480 44312 5442
rect 47596 4146 47624 147018
rect 50344 145920 50396 145926
rect 50344 145862 50396 145868
rect 47860 7608 47912 7614
rect 47860 7550 47912 7556
rect 45468 4140 45520 4146
rect 45468 4082 45520 4088
rect 47584 4140 47636 4146
rect 47584 4082 47636 4088
rect 45480 480 45508 4082
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 46676 480 46704 3878
rect 47872 480 47900 7550
rect 48964 6180 49016 6186
rect 48964 6122 49016 6128
rect 48976 480 49004 6122
rect 50356 4010 50384 145862
rect 50344 4004 50396 4010
rect 50344 3946 50396 3952
rect 52380 3398 52408 147154
rect 53104 145852 53156 145858
rect 53104 145794 53156 145800
rect 52552 6248 52604 6254
rect 52552 6190 52604 6196
rect 51356 3392 51408 3398
rect 51356 3334 51408 3340
rect 52368 3392 52420 3398
rect 52368 3334 52420 3340
rect 50160 2984 50212 2990
rect 50160 2926 50212 2932
rect 50172 480 50200 2926
rect 51368 480 51396 3334
rect 52564 480 52592 6190
rect 53116 2990 53144 145794
rect 57244 144220 57296 144226
rect 57244 144162 57296 144168
rect 54944 10328 54996 10334
rect 54944 10270 54996 10276
rect 53748 3188 53800 3194
rect 53748 3130 53800 3136
rect 53104 2984 53156 2990
rect 53104 2926 53156 2932
rect 53760 480 53788 3130
rect 54956 480 54984 10270
rect 57256 6914 57284 144162
rect 57164 6886 57284 6914
rect 56048 6316 56100 6322
rect 56048 6258 56100 6264
rect 56060 480 56088 6258
rect 57164 3194 57192 6886
rect 57244 4004 57296 4010
rect 57244 3946 57296 3952
rect 57152 3188 57204 3194
rect 57152 3130 57204 3136
rect 57256 480 57284 3946
rect 59280 3398 59308 147290
rect 62028 147280 62080 147286
rect 62028 147222 62080 147228
rect 60832 8968 60884 8974
rect 60832 8910 60884 8916
rect 59636 6384 59688 6390
rect 59636 6326 59688 6332
rect 58440 3392 58492 3398
rect 58440 3334 58492 3340
rect 59268 3392 59320 3398
rect 59268 3334 59320 3340
rect 58452 480 58480 3334
rect 59648 480 59676 6326
rect 60844 480 60872 8910
rect 62040 480 62068 147222
rect 65524 146056 65576 146062
rect 65524 145998 65576 146004
rect 65536 6914 65564 145998
rect 71044 145988 71096 145994
rect 71044 145930 71096 145936
rect 68284 144288 68336 144294
rect 68284 144230 68336 144236
rect 65444 6886 65564 6914
rect 63224 6452 63276 6458
rect 63224 6394 63276 6400
rect 63236 480 63264 6394
rect 64328 4072 64380 4078
rect 64328 4014 64380 4020
rect 64340 480 64368 4014
rect 65444 4010 65472 6886
rect 66720 6520 66772 6526
rect 66720 6462 66772 6468
rect 65524 4752 65576 4758
rect 65524 4694 65576 4700
rect 65432 4004 65484 4010
rect 65432 3946 65484 3952
rect 65536 480 65564 4694
rect 66732 480 66760 6462
rect 68296 4078 68324 144230
rect 70308 6588 70360 6594
rect 70308 6530 70360 6536
rect 69112 4548 69164 4554
rect 69112 4490 69164 4496
rect 68284 4072 68336 4078
rect 68284 4014 68336 4020
rect 67916 3392 67968 3398
rect 67916 3334 67968 3340
rect 67928 480 67956 3334
rect 69124 480 69152 4490
rect 70320 480 70348 6530
rect 71056 3398 71084 145930
rect 72424 144356 72476 144362
rect 72424 144298 72476 144304
rect 72436 3398 72464 144298
rect 75196 4690 75224 148786
rect 88248 147416 88300 147422
rect 88248 147358 88300 147364
rect 76564 146124 76616 146130
rect 76564 146066 76616 146072
rect 73804 4684 73856 4690
rect 73804 4626 73856 4632
rect 75184 4684 75236 4690
rect 75184 4626 75236 4632
rect 72608 4616 72660 4622
rect 72608 4558 72660 4564
rect 71044 3392 71096 3398
rect 71044 3334 71096 3340
rect 71504 3392 71556 3398
rect 71504 3334 71556 3340
rect 72424 3392 72476 3398
rect 72424 3334 72476 3340
rect 71516 480 71544 3334
rect 72620 480 72648 4558
rect 73816 480 73844 4626
rect 76196 4480 76248 4486
rect 76196 4422 76248 4428
rect 75000 3392 75052 3398
rect 75000 3334 75052 3340
rect 75012 480 75040 3334
rect 76208 480 76236 4422
rect 76576 3398 76604 146066
rect 80888 7676 80940 7682
rect 80888 7618 80940 7624
rect 77392 6656 77444 6662
rect 77392 6598 77444 6604
rect 76564 3392 76616 3398
rect 76564 3334 76616 3340
rect 77404 480 77432 6598
rect 79692 4480 79744 4486
rect 79692 4422 79744 4428
rect 78588 4004 78640 4010
rect 78588 3946 78640 3952
rect 78600 480 78628 3946
rect 79704 480 79732 4422
rect 80900 480 80928 7618
rect 88260 6914 88288 147358
rect 87984 6886 88288 6914
rect 84476 6724 84528 6730
rect 84476 6666 84528 6672
rect 83280 4412 83332 4418
rect 83280 4354 83332 4360
rect 82084 4072 82136 4078
rect 82084 4014 82136 4020
rect 82096 480 82124 4014
rect 83292 480 83320 4354
rect 84488 480 84516 6666
rect 86868 4344 86920 4350
rect 86868 4286 86920 4292
rect 85672 3392 85724 3398
rect 85672 3334 85724 3340
rect 85684 480 85712 3334
rect 86880 480 86908 4286
rect 87984 480 88012 6886
rect 93136 5574 93164 148854
rect 99288 147552 99340 147558
rect 99288 147494 99340 147500
rect 95148 147484 95200 147490
rect 95148 147426 95200 147432
rect 95056 9036 95108 9042
rect 95056 8978 95108 8984
rect 91560 5568 91612 5574
rect 91560 5510 91612 5516
rect 93124 5568 93176 5574
rect 93124 5510 93176 5516
rect 90364 4276 90416 4282
rect 90364 4218 90416 4224
rect 89168 3256 89220 3262
rect 89168 3198 89220 3204
rect 89180 480 89208 3198
rect 90376 480 90404 4218
rect 91572 480 91600 5510
rect 93952 4140 94004 4146
rect 93952 4082 94004 4088
rect 92756 3324 92808 3330
rect 92756 3266 92808 3272
rect 92768 480 92796 3266
rect 93964 480 93992 4082
rect 95068 3482 95096 8978
rect 95160 4146 95188 147426
rect 97448 6792 97500 6798
rect 97448 6734 97500 6740
rect 95148 4140 95200 4146
rect 95148 4082 95200 4088
rect 95068 3454 95188 3482
rect 95160 480 95188 3454
rect 96252 3188 96304 3194
rect 96252 3130 96304 3136
rect 96264 480 96292 3130
rect 97460 480 97488 6734
rect 99300 3262 99328 147494
rect 101036 6112 101088 6118
rect 101036 6054 101088 6060
rect 98644 3256 98696 3262
rect 98644 3198 98696 3204
rect 99288 3256 99340 3262
rect 99288 3198 99340 3204
rect 98656 480 98684 3198
rect 99840 3188 99892 3194
rect 99840 3130 99892 3136
rect 99852 480 99880 3130
rect 101048 480 101076 6054
rect 104176 5574 104204 148922
rect 106188 147620 106240 147626
rect 106188 147562 106240 147568
rect 104532 6044 104584 6050
rect 104532 5986 104584 5992
rect 102232 5568 102284 5574
rect 102232 5510 102284 5516
rect 104164 5568 104216 5574
rect 104164 5510 104216 5516
rect 102244 480 102272 5510
rect 103336 3120 103388 3126
rect 103336 3062 103388 3068
rect 103348 480 103376 3062
rect 104544 480 104572 5986
rect 106200 3058 106228 147562
rect 107580 3058 107608 148990
rect 111064 148300 111116 148306
rect 111064 148242 111116 148248
rect 108120 5976 108172 5982
rect 108120 5918 108172 5924
rect 105728 3052 105780 3058
rect 105728 2994 105780 3000
rect 106188 3052 106240 3058
rect 106188 2994 106240 3000
rect 106924 3052 106976 3058
rect 106924 2994 106976 3000
rect 107568 3052 107620 3058
rect 107568 2994 107620 3000
rect 105740 480 105768 2994
rect 106936 480 106964 2994
rect 108132 480 108160 5918
rect 111076 5574 111104 148242
rect 114468 148232 114520 148238
rect 114468 148174 114520 148180
rect 113088 146872 113140 146878
rect 113088 146814 113140 146820
rect 113100 6914 113128 146814
rect 112824 6886 113128 6914
rect 111616 5908 111668 5914
rect 111616 5850 111668 5856
rect 109316 5568 109368 5574
rect 109316 5510 109368 5516
rect 111064 5568 111116 5574
rect 111064 5510 111116 5516
rect 109328 480 109356 5510
rect 110512 3052 110564 3058
rect 110512 2994 110564 3000
rect 110524 480 110552 2994
rect 111628 480 111656 5850
rect 112824 480 112852 6886
rect 114480 2990 114508 148174
rect 115204 148096 115256 148102
rect 115204 148038 115256 148044
rect 115216 7682 115244 148038
rect 116584 148028 116636 148034
rect 116584 147970 116636 147976
rect 116596 10334 116624 147970
rect 119356 137970 119384 557806
rect 122116 346390 122144 559370
rect 155132 559156 155184 559162
rect 155132 559098 155184 559104
rect 123484 558068 123536 558074
rect 123484 558010 123536 558016
rect 122104 346384 122156 346390
rect 122104 346326 122156 346332
rect 123496 241466 123524 558010
rect 155144 557940 155172 559098
rect 167012 557940 167040 560594
rect 172980 559224 173032 559230
rect 172980 559166 173032 559172
rect 169944 559020 169996 559026
rect 169944 558962 169996 558968
rect 169956 557940 169984 558962
rect 172992 557940 173020 559166
rect 175936 557940 175964 560662
rect 178868 558136 178920 558142
rect 178868 558078 178920 558084
rect 178880 557940 178908 558078
rect 184860 557940 184888 560730
rect 190736 559360 190788 559366
rect 190736 559302 190788 559308
rect 187792 558204 187844 558210
rect 187792 558146 187844 558152
rect 187804 557940 187832 558146
rect 190748 557940 190776 559302
rect 193692 557940 193720 560798
rect 196716 559496 196768 559502
rect 196716 559438 196768 559444
rect 196728 557940 196756 559438
rect 199844 558000 199896 558006
rect 199686 557948 199844 557954
rect 199686 557942 199896 557948
rect 199686 557926 199884 557942
rect 202616 557940 202644 560866
rect 205548 559632 205600 559638
rect 205548 559574 205600 559580
rect 205560 557940 205588 559574
rect 211540 557940 211568 561002
rect 214472 558272 214524 558278
rect 214472 558214 214524 558220
rect 214484 557940 214512 558214
rect 232332 557940 232360 563042
rect 235736 557954 235764 567166
rect 235920 561474 235948 699654
rect 253848 696992 253900 696998
rect 253848 696934 253900 696940
rect 251088 670812 251140 670818
rect 251088 670754 251140 670760
rect 244188 643136 244240 643142
rect 244188 643078 244240 643084
rect 241428 616888 241480 616894
rect 241428 616830 241480 616836
rect 238668 576904 238720 576910
rect 238668 576846 238720 576852
rect 235908 561468 235960 561474
rect 235908 561410 235960 561416
rect 238680 557954 238708 576846
rect 241440 557954 241468 616830
rect 235290 557926 235764 557954
rect 238234 557926 238708 557954
rect 241178 557926 241468 557954
rect 244200 557940 244228 643078
rect 248328 630692 248380 630698
rect 248328 630634 248380 630640
rect 248340 561678 248368 630634
rect 251100 561678 251128 670754
rect 253860 561678 253888 696934
rect 256608 683256 256660 683262
rect 256608 683198 256660 683204
rect 256620 567194 256648 683198
rect 256528 567166 256648 567194
rect 247132 561672 247184 561678
rect 247132 561614 247184 561620
rect 248328 561672 248380 561678
rect 248328 561614 248380 561620
rect 250076 561672 250128 561678
rect 250076 561614 250128 561620
rect 251088 561672 251140 561678
rect 251088 561614 251140 561620
rect 253020 561672 253072 561678
rect 253020 561614 253072 561620
rect 253848 561672 253900 561678
rect 253848 561614 253900 561620
rect 247144 557940 247172 561614
rect 250088 557940 250116 561614
rect 253032 557940 253060 561614
rect 256528 557954 256556 567166
rect 259000 560992 259052 560998
rect 259000 560934 259052 560940
rect 256082 557926 256556 557954
rect 259012 557940 259040 560934
rect 262140 557954 262168 700538
rect 264888 700528 264940 700534
rect 264888 700470 264940 700476
rect 261970 557926 262168 557954
rect 264900 557940 264928 700470
rect 267660 699854 267688 703520
rect 271788 700868 271840 700874
rect 271788 700810 271840 700816
rect 267648 699848 267700 699854
rect 267648 699790 267700 699796
rect 271800 561678 271828 700810
rect 274548 700800 274600 700806
rect 274548 700742 274600 700748
rect 274560 561678 274588 700742
rect 282828 700256 282880 700262
rect 282828 700198 282880 700204
rect 280068 700188 280120 700194
rect 280068 700130 280120 700136
rect 270868 561672 270920 561678
rect 270868 561614 270920 561620
rect 271788 561672 271840 561678
rect 271788 561614 271840 561620
rect 273812 561672 273864 561678
rect 273812 561614 273864 561620
rect 274548 561672 274600 561678
rect 274548 561614 274600 561620
rect 267924 561128 267976 561134
rect 267924 561070 267976 561076
rect 267936 557940 267964 561070
rect 270880 557940 270908 561614
rect 273824 557940 273852 561614
rect 276756 561264 276808 561270
rect 276756 561206 276808 561212
rect 276768 557940 276796 561206
rect 280080 557954 280108 700130
rect 282840 557954 282868 700198
rect 283852 699786 283880 703520
rect 292488 699984 292540 699990
rect 292488 699926 292540 699932
rect 289728 699916 289780 699922
rect 289728 699858 289780 699864
rect 283840 699780 283892 699786
rect 283840 699722 283892 699728
rect 289740 561678 289768 699858
rect 292500 561678 292528 699926
rect 296720 699848 296772 699854
rect 296720 699790 296772 699796
rect 296732 576854 296760 699790
rect 296732 576826 297128 576854
rect 288624 561672 288676 561678
rect 288624 561614 288676 561620
rect 289728 561672 289780 561678
rect 289728 561614 289780 561620
rect 291660 561672 291712 561678
rect 291660 561614 291712 561620
rect 292488 561672 292540 561678
rect 292488 561614 292540 561620
rect 285680 561400 285732 561406
rect 285680 561342 285732 561348
rect 279818 557926 280108 557954
rect 282762 557926 282868 557954
rect 285692 557940 285720 561342
rect 288636 557940 288664 561614
rect 291672 557940 291700 561614
rect 294604 561536 294656 561542
rect 294604 561478 294656 561484
rect 294616 557940 294644 561478
rect 297100 557954 297128 576826
rect 299492 561542 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 317420 701004 317472 701010
rect 317420 700946 317472 700952
rect 314660 700936 314712 700942
rect 314660 700878 314712 700884
rect 306380 700120 306432 700126
rect 306380 700062 306432 700068
rect 299572 699780 299624 699786
rect 299572 699722 299624 699728
rect 299584 576854 299612 699722
rect 299584 576826 300256 576854
rect 299480 561536 299532 561542
rect 299480 561478 299532 561484
rect 300228 557954 300256 576826
rect 303528 561468 303580 561474
rect 303528 561410 303580 561416
rect 297100 557926 297574 557954
rect 300228 557926 300610 557954
rect 303540 557940 303568 561410
rect 306392 557954 306420 700062
rect 309140 700052 309192 700058
rect 309140 699994 309192 700000
rect 309152 557954 309180 699994
rect 314672 576854 314700 700878
rect 317432 576854 317460 700946
rect 327080 700732 327132 700738
rect 327080 700674 327132 700680
rect 324320 700664 324372 700670
rect 324320 700606 324372 700612
rect 314672 576826 314976 576854
rect 317432 576826 317920 576854
rect 312452 561332 312504 561338
rect 312452 561274 312504 561280
rect 306392 557926 306498 557954
rect 309152 557926 309442 557954
rect 312464 557940 312492 561274
rect 314948 557954 314976 576826
rect 317892 557954 317920 576826
rect 321284 561196 321336 561202
rect 321284 561138 321336 561144
rect 314948 557926 315422 557954
rect 317892 557926 318366 557954
rect 321296 557940 321324 561138
rect 324332 557940 324360 700606
rect 327092 557954 327120 700674
rect 329840 700460 329892 700466
rect 329840 700402 329892 700408
rect 329852 557954 329880 700402
rect 332520 699922 332548 703520
rect 335360 700392 335412 700398
rect 335360 700334 335412 700340
rect 332600 700324 332652 700330
rect 332600 700266 332652 700272
rect 332508 699916 332560 699922
rect 332508 699858 332560 699864
rect 332612 576854 332640 700266
rect 335372 576854 335400 700334
rect 348804 699990 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 699984 348844 699990
rect 348792 699926 348844 699932
rect 338120 683188 338172 683194
rect 338120 683130 338172 683136
rect 338132 576854 338160 683130
rect 345020 670744 345072 670750
rect 345020 670686 345072 670692
rect 340880 656940 340932 656946
rect 340880 656882 340932 656888
rect 340892 576854 340920 656882
rect 332612 576826 332824 576854
rect 335372 576826 335768 576854
rect 338132 576826 338712 576854
rect 340892 576826 341656 576854
rect 332796 557954 332824 576826
rect 335740 557954 335768 576826
rect 338684 557954 338712 576826
rect 341628 557954 341656 576826
rect 327092 557926 327290 557954
rect 329852 557926 330234 557954
rect 332796 557926 333178 557954
rect 335740 557926 336214 557954
rect 338684 557926 339158 557954
rect 341628 557926 342102 557954
rect 345032 557940 345060 670686
rect 347780 632120 347832 632126
rect 347780 632062 347832 632068
rect 347792 557954 347820 632062
rect 353300 618316 353352 618322
rect 353300 618258 353352 618264
rect 350540 605872 350592 605878
rect 350540 605814 350592 605820
rect 350552 576854 350580 605814
rect 353312 576854 353340 618258
rect 356060 579692 356112 579698
rect 356060 579634 356112 579640
rect 356072 576854 356100 579634
rect 350552 576826 350672 576854
rect 353312 576826 353616 576854
rect 356072 576826 356560 576854
rect 350644 557954 350672 576826
rect 353588 557954 353616 576826
rect 356532 557954 356560 576826
rect 362868 565888 362920 565894
rect 362868 565830 362920 565836
rect 347792 557926 348082 557954
rect 350644 557926 351026 557954
rect 353588 557926 353970 557954
rect 356532 557926 356914 557954
rect 362880 557940 362908 565830
rect 364352 561406 364380 702406
rect 397472 700194 397500 703520
rect 413664 700262 413692 703520
rect 413652 700256 413704 700262
rect 413652 700198 413704 700204
rect 397460 700188 397512 700194
rect 397460 700130 397512 700136
rect 364340 561400 364392 561406
rect 364340 561342 364392 561348
rect 429212 561270 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 700874 462360 703520
rect 462320 700868 462372 700874
rect 462320 700810 462372 700816
rect 478524 700806 478552 703520
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 429200 561264 429252 561270
rect 429200 561206 429252 561212
rect 494072 561134 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 700602 527220 703520
rect 527180 700596 527232 700602
rect 527180 700538 527232 700544
rect 543476 700534 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700528 543516 700534
rect 543464 700470 543516 700476
rect 494060 561128 494112 561134
rect 494060 561070 494112 561076
rect 486424 561060 486476 561066
rect 486424 561002 486476 561008
rect 485044 560924 485096 560930
rect 485044 560866 485096 560872
rect 483664 560856 483716 560862
rect 483664 560798 483716 560804
rect 482284 560788 482336 560794
rect 482284 560730 482336 560736
rect 479524 560720 479576 560726
rect 479524 560662 479576 560668
rect 475384 560652 475436 560658
rect 475384 560594 475436 560600
rect 398472 560584 398524 560590
rect 398472 560526 398524 560532
rect 380624 559564 380676 559570
rect 380624 559506 380676 559512
rect 380636 557940 380664 559506
rect 395528 559428 395580 559434
rect 395528 559370 395580 559376
rect 386432 557938 386630 557954
rect 395540 557940 395568 559370
rect 398484 557940 398512 560526
rect 407396 560516 407448 560522
rect 407396 560458 407448 560464
rect 407408 557940 407436 560458
rect 416228 560448 416280 560454
rect 416228 560390 416280 560396
rect 410340 558952 410392 558958
rect 410340 558894 410392 558900
rect 410352 557940 410380 558894
rect 412916 558068 412968 558074
rect 412916 558010 412968 558016
rect 412928 557954 412956 558010
rect 386420 557932 386630 557938
rect 386472 557926 386630 557932
rect 412928 557926 413310 557954
rect 416240 557940 416268 560390
rect 425152 560380 425204 560386
rect 425152 560322 425204 560328
rect 422208 559292 422260 559298
rect 422208 559234 422260 559240
rect 422220 557940 422248 559234
rect 425164 557940 425192 560322
rect 434076 560312 434128 560318
rect 434076 560254 434128 560260
rect 428096 559088 428148 559094
rect 428096 559030 428148 559036
rect 428108 557940 428136 559030
rect 434088 557940 434116 560254
rect 468484 559632 468536 559638
rect 468484 559574 468536 559580
rect 467104 559496 467156 559502
rect 467104 559438 467156 559444
rect 462964 558272 463016 558278
rect 462964 558214 463016 558220
rect 386420 557874 386472 557880
rect 430764 557864 430816 557870
rect 181838 557802 182128 557818
rect 430816 557812 431158 557818
rect 430764 557806 431158 557812
rect 181838 557796 182140 557802
rect 181838 557790 182088 557796
rect 430776 557790 431158 557806
rect 182088 557738 182140 557744
rect 164148 557728 164200 557734
rect 128478 557666 128768 557682
rect 164082 557676 164148 557682
rect 164082 557670 164200 557676
rect 128478 557660 128780 557666
rect 128478 557654 128728 557660
rect 164082 557654 164188 557670
rect 128728 557602 128780 557608
rect 418988 557592 419040 557598
rect 131670 557560 131726 557569
rect 131422 557518 131670 557546
rect 134614 557560 134670 557569
rect 134366 557518 134614 557546
rect 131670 557495 131726 557504
rect 137742 557560 137798 557569
rect 137402 557518 137742 557546
rect 134614 557495 134670 557504
rect 140594 557560 140650 557569
rect 140346 557518 140594 557546
rect 137742 557495 137798 557504
rect 143354 557560 143410 557569
rect 143290 557518 143354 557546
rect 140594 557495 140650 557504
rect 143354 557495 143410 557504
rect 145930 557560 145986 557569
rect 149334 557560 149390 557569
rect 145986 557518 146234 557546
rect 149270 557518 149334 557546
rect 145930 557495 145986 557504
rect 152462 557560 152518 557569
rect 152214 557518 152462 557546
rect 149334 557495 149390 557504
rect 158350 557560 158406 557569
rect 158102 557518 158350 557546
rect 152462 557495 152518 557504
rect 436650 557560 436706 557569
rect 419040 557540 419290 557546
rect 418988 557534 419290 557540
rect 419000 557518 419290 557534
rect 158350 557495 158406 557504
rect 439594 557560 439650 557569
rect 436706 557518 437046 557546
rect 436650 557495 436706 557504
rect 443090 557560 443146 557569
rect 439650 557518 439990 557546
rect 443026 557518 443090 557546
rect 439594 557495 439650 557504
rect 443090 557495 443146 557504
rect 445758 557560 445814 557569
rect 448610 557560 448666 557569
rect 445814 557518 445970 557546
rect 445758 557495 445814 557504
rect 451554 557560 451610 557569
rect 448666 557518 448914 557546
rect 448610 557495 448666 557504
rect 454498 557560 454554 557569
rect 451610 557518 451858 557546
rect 451554 557495 451610 557504
rect 457442 557560 457498 557569
rect 454554 557518 454894 557546
rect 454498 557495 454554 557504
rect 460386 557560 460442 557569
rect 457498 557518 457838 557546
rect 457442 557495 457498 557504
rect 460442 557518 460782 557546
rect 460386 557495 460442 557504
rect 359556 557456 359608 557462
rect 124232 557382 125534 557410
rect 161138 557394 161336 557410
rect 208610 557394 208992 557410
rect 217442 557394 217824 557410
rect 220478 557394 220768 557410
rect 223422 557394 223528 557410
rect 226366 557394 226656 557410
rect 229310 557394 229600 557410
rect 365628 557456 365680 557462
rect 359608 557404 359950 557410
rect 359556 557398 359950 557404
rect 368480 557456 368532 557462
rect 365680 557404 365838 557410
rect 365628 557398 365838 557404
rect 371516 557456 371568 557462
rect 368532 557404 368782 557410
rect 368480 557398 368782 557404
rect 374460 557456 374512 557462
rect 371568 557404 371818 557410
rect 371516 557398 371818 557404
rect 377404 557456 377456 557462
rect 374512 557404 374762 557410
rect 374460 557398 374762 557404
rect 383752 557456 383804 557462
rect 377456 557404 377706 557410
rect 377404 557398 377706 557404
rect 161138 557388 161348 557394
rect 161138 557382 161296 557388
rect 123484 241460 123536 241466
rect 123484 241402 123536 241408
rect 119436 148164 119488 148170
rect 119436 148106 119488 148112
rect 119344 137964 119396 137970
rect 119344 137906 119396 137912
rect 116584 10328 116636 10334
rect 116584 10270 116636 10276
rect 119448 8294 119476 148106
rect 122104 147960 122156 147966
rect 122104 147902 122156 147908
rect 119988 141432 120040 141438
rect 119988 141374 120040 141380
rect 116400 8288 116452 8294
rect 116400 8230 116452 8236
rect 119436 8288 119488 8294
rect 119436 8230 119488 8236
rect 115204 7676 115256 7682
rect 115204 7618 115256 7624
rect 115204 5840 115256 5846
rect 115204 5782 115256 5788
rect 114008 2984 114060 2990
rect 114008 2926 114060 2932
rect 114468 2984 114520 2990
rect 114468 2926 114520 2932
rect 114020 480 114048 2926
rect 115216 480 115244 5782
rect 116412 480 116440 8230
rect 120000 6914 120028 141374
rect 122116 7614 122144 147902
rect 123484 147688 123536 147694
rect 123484 147630 123536 147636
rect 123496 91798 123524 147630
rect 124128 146192 124180 146198
rect 124128 146134 124180 146140
rect 123484 91792 123536 91798
rect 123484 91734 123536 91740
rect 122104 7608 122156 7614
rect 122104 7550 122156 7556
rect 119908 6886 120028 6914
rect 118792 5772 118844 5778
rect 118792 5714 118844 5720
rect 117596 2848 117648 2854
rect 117596 2790 117648 2796
rect 117608 480 117636 2790
rect 118804 480 118832 5714
rect 119908 480 119936 6886
rect 122288 5704 122340 5710
rect 122288 5646 122340 5652
rect 121092 2916 121144 2922
rect 121092 2858 121144 2864
rect 121104 480 121132 2858
rect 122300 480 122328 5646
rect 124140 2990 124168 146134
rect 124232 6866 124260 557382
rect 208610 557388 209004 557394
rect 208610 557382 208952 557388
rect 161296 557330 161348 557336
rect 217442 557388 217836 557394
rect 217442 557382 217784 557388
rect 208952 557330 209004 557336
rect 220478 557388 220780 557394
rect 220478 557382 220728 557388
rect 217784 557330 217836 557336
rect 223422 557388 223540 557394
rect 223422 557382 223488 557388
rect 220728 557330 220780 557336
rect 226366 557388 226668 557394
rect 226366 557382 226616 557388
rect 223488 557330 223540 557336
rect 229310 557388 229612 557394
rect 229310 557382 229560 557388
rect 226616 557330 226668 557336
rect 359568 557382 359950 557398
rect 365640 557382 365838 557398
rect 368492 557382 368782 557398
rect 371528 557382 371818 557398
rect 374472 557382 374762 557398
rect 377416 557382 377706 557398
rect 383686 557404 383752 557410
rect 383686 557398 383804 557404
rect 389180 557456 389232 557462
rect 392124 557456 392176 557462
rect 389232 557404 389574 557410
rect 389180 557398 389574 557404
rect 401140 557456 401192 557462
rect 392176 557404 392518 557410
rect 392124 557398 392518 557404
rect 404176 557456 404228 557462
rect 401192 557404 401442 557410
rect 401140 557398 401442 557404
rect 404228 557404 404386 557410
rect 404176 557398 404386 557404
rect 383686 557382 383792 557398
rect 389192 557382 389574 557398
rect 392136 557382 392518 557398
rect 401152 557382 401442 557398
rect 404188 557382 404386 557398
rect 229560 557330 229612 557336
rect 462976 458182 463004 558214
rect 465724 558204 465776 558210
rect 465724 558146 465776 558152
rect 464344 558136 464396 558142
rect 464344 558078 464396 558084
rect 462964 458176 463016 458182
rect 462964 458118 463016 458124
rect 464356 245614 464384 558078
rect 465736 299470 465764 558146
rect 467116 353258 467144 559438
rect 468496 405686 468524 559574
rect 472624 559156 472676 559162
rect 472624 559098 472676 559104
rect 471244 557660 471296 557666
rect 471244 557602 471296 557608
rect 468484 405680 468536 405686
rect 468484 405622 468536 405628
rect 467104 353252 467156 353258
rect 467104 353194 467156 353200
rect 465724 299464 465776 299470
rect 465724 299406 465776 299412
rect 464344 245608 464396 245614
rect 464344 245550 464396 245556
rect 124324 148578 124352 150484
rect 124968 148714 124996 150484
rect 124956 148708 125008 148714
rect 124956 148650 125008 148656
rect 124312 148572 124364 148578
rect 124312 148514 124364 148520
rect 125612 147694 125640 150484
rect 125704 150470 126362 150498
rect 127006 150470 127204 150498
rect 125600 147688 125652 147694
rect 125600 147630 125652 147636
rect 124220 6860 124272 6866
rect 124220 6802 124272 6808
rect 125704 4826 125732 150470
rect 126980 7676 127032 7682
rect 126980 7618 127032 7624
rect 125876 7608 125928 7614
rect 125876 7550 125928 7556
rect 125692 4820 125744 4826
rect 125692 4762 125744 4768
rect 123484 2984 123536 2990
rect 123484 2926 123536 2932
rect 124128 2984 124180 2990
rect 124128 2926 124180 2932
rect 123496 480 123524 2926
rect 124680 2780 124732 2786
rect 124680 2722 124732 2728
rect 124692 480 124720 2722
rect 125888 480 125916 7550
rect 126992 480 127020 7618
rect 127176 3369 127204 150470
rect 127728 148374 127756 150484
rect 128372 148442 128400 150484
rect 128464 150470 129122 150498
rect 128360 148436 128412 148442
rect 128360 148378 128412 148384
rect 127716 148368 127768 148374
rect 127716 148310 127768 148316
rect 128464 4894 128492 150470
rect 129004 148368 129056 148374
rect 129004 148310 129056 148316
rect 128452 4888 128504 4894
rect 128452 4830 128504 4836
rect 129016 4214 129044 148310
rect 129752 145586 129780 150484
rect 129936 150470 130502 150498
rect 131146 150470 131252 150498
rect 129740 145580 129792 145586
rect 129740 145522 129792 145528
rect 129372 6928 129424 6934
rect 129372 6870 129424 6876
rect 128176 4208 128228 4214
rect 128176 4150 128228 4156
rect 129004 4208 129056 4214
rect 129004 4150 129056 4156
rect 127162 3360 127218 3369
rect 127162 3295 127218 3304
rect 128188 480 128216 4150
rect 129384 480 129412 6870
rect 129936 3505 129964 150470
rect 130568 7744 130620 7750
rect 130568 7686 130620 7692
rect 129922 3496 129978 3505
rect 129922 3431 129978 3440
rect 130580 480 130608 7686
rect 131224 4962 131252 150470
rect 131868 148646 131896 150484
rect 132526 150470 132632 150498
rect 131856 148640 131908 148646
rect 131856 148582 131908 148588
rect 131212 4956 131264 4962
rect 131212 4898 131264 4904
rect 131764 4888 131816 4894
rect 131764 4830 131816 4836
rect 131776 480 131804 4830
rect 132604 3641 132632 150470
rect 133156 148510 133184 150484
rect 133906 150470 134012 150498
rect 133144 148504 133196 148510
rect 133144 148446 133196 148452
rect 133328 148504 133380 148510
rect 133328 148446 133380 148452
rect 133236 148436 133288 148442
rect 133236 148378 133288 148384
rect 133248 145330 133276 148378
rect 133156 145302 133276 145330
rect 133156 4894 133184 145302
rect 133340 142154 133368 148446
rect 133248 142126 133368 142154
rect 133248 6934 133276 142126
rect 133420 11756 133472 11762
rect 133420 11698 133472 11704
rect 133236 6928 133288 6934
rect 133236 6870 133288 6876
rect 133144 4888 133196 4894
rect 133144 4830 133196 4836
rect 132590 3632 132646 3641
rect 132590 3567 132646 3576
rect 132972 598 133184 626
rect 132972 480 133000 598
rect 133156 490 133184 598
rect 133432 490 133460 11698
rect 133984 4826 134012 150470
rect 134536 146946 134564 150484
rect 135272 148782 135300 150484
rect 135364 150470 135930 150498
rect 135260 148776 135312 148782
rect 135260 148718 135312 148724
rect 134524 146940 134576 146946
rect 134524 146882 134576 146888
rect 135260 7880 135312 7886
rect 135260 7822 135312 7828
rect 134156 7812 134208 7818
rect 134156 7754 134208 7760
rect 133972 4820 134024 4826
rect 133972 4762 134024 4768
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133156 462 133460 490
rect 134168 480 134196 7754
rect 135272 480 135300 7822
rect 135364 3777 135392 150470
rect 136652 5098 136680 150484
rect 137296 145722 137324 150484
rect 137284 145716 137336 145722
rect 137284 145658 137336 145664
rect 138032 142186 138060 150484
rect 138124 150470 138690 150498
rect 139426 150470 139532 150498
rect 138020 142180 138072 142186
rect 138020 142122 138072 142128
rect 137652 15904 137704 15910
rect 137652 15846 137704 15852
rect 136640 5092 136692 5098
rect 136640 5034 136692 5040
rect 136456 4888 136508 4894
rect 136456 4830 136508 4836
rect 135350 3768 135406 3777
rect 135350 3703 135406 3712
rect 136468 480 136496 4830
rect 137664 480 137692 15846
rect 138124 3534 138152 150470
rect 138204 142180 138256 142186
rect 138204 142122 138256 142128
rect 138112 3528 138164 3534
rect 138112 3470 138164 3476
rect 138216 3466 138244 142122
rect 138848 8016 138900 8022
rect 138848 7958 138900 7964
rect 138204 3460 138256 3466
rect 138204 3402 138256 3408
rect 138860 480 138888 7958
rect 139504 5166 139532 150470
rect 140056 147014 140084 150484
rect 140044 147008 140096 147014
rect 140044 146950 140096 146956
rect 140792 142186 140820 150484
rect 140884 150470 141450 150498
rect 140780 142180 140832 142186
rect 140780 142122 140832 142128
rect 140044 7948 140096 7954
rect 140044 7890 140096 7896
rect 139492 5160 139544 5166
rect 139492 5102 139544 5108
rect 140056 480 140084 7890
rect 140884 5234 140912 150470
rect 142080 145654 142108 150484
rect 142172 150470 142830 150498
rect 142908 150470 143474 150498
rect 142068 145648 142120 145654
rect 142068 145590 142120 145596
rect 140964 142180 141016 142186
rect 140964 142122 141016 142128
rect 140872 5228 140924 5234
rect 140872 5170 140924 5176
rect 140976 3602 141004 142122
rect 141240 4820 141292 4826
rect 141240 4762 141292 4768
rect 140964 3596 141016 3602
rect 140964 3538 141016 3544
rect 141252 480 141280 4762
rect 142172 3670 142200 150470
rect 142908 142154 142936 150470
rect 144196 145790 144224 150484
rect 144288 150470 144854 150498
rect 145024 150470 145590 150498
rect 144184 145784 144236 145790
rect 144184 145726 144236 145732
rect 144288 145636 144316 150470
rect 144368 148640 144420 148646
rect 144368 148582 144420 148588
rect 142264 142126 142936 142154
rect 143552 145608 144316 145636
rect 142264 5302 142292 142126
rect 143552 16574 143580 145608
rect 144380 142154 144408 148582
rect 144196 142126 144408 142154
rect 143552 16546 143672 16574
rect 142436 9172 142488 9178
rect 142436 9114 142488 9120
rect 142252 5296 142304 5302
rect 142252 5238 142304 5244
rect 142160 3664 142212 3670
rect 142160 3606 142212 3612
rect 142448 480 142476 9114
rect 143540 4208 143592 4214
rect 143540 4150 143592 4156
rect 143552 480 143580 4150
rect 143644 3806 143672 16546
rect 144196 4894 144224 142126
rect 145024 5370 145052 150470
rect 146220 147150 146248 150484
rect 146312 150470 146970 150498
rect 147048 150470 147614 150498
rect 146208 147144 146260 147150
rect 146208 147086 146260 147092
rect 145932 9104 145984 9110
rect 145932 9046 145984 9052
rect 145012 5364 145064 5370
rect 145012 5306 145064 5312
rect 144184 4888 144236 4894
rect 144184 4830 144236 4836
rect 144736 4888 144788 4894
rect 144736 4830 144788 4836
rect 143632 3800 143684 3806
rect 143632 3742 143684 3748
rect 144748 480 144776 4830
rect 145944 480 145972 9046
rect 146312 3738 146340 150470
rect 147048 146418 147076 150470
rect 147128 148572 147180 148578
rect 147128 148514 147180 148520
rect 146404 146390 147076 146418
rect 146404 5438 146432 146390
rect 147140 142154 147168 148514
rect 148336 145926 148364 150484
rect 148428 150470 148994 150498
rect 149164 150470 149638 150498
rect 148324 145920 148376 145926
rect 148324 145862 148376 145868
rect 148428 142154 148456 150470
rect 146956 142126 147168 142154
rect 147692 142126 148456 142154
rect 146392 5432 146444 5438
rect 146392 5374 146444 5380
rect 146956 4214 146984 142126
rect 147128 8084 147180 8090
rect 147128 8026 147180 8032
rect 146944 4208 146996 4214
rect 146944 4150 146996 4156
rect 146300 3732 146352 3738
rect 146300 3674 146352 3680
rect 147140 480 147168 8026
rect 147692 3874 147720 142126
rect 149164 5506 149192 150470
rect 150360 147082 150388 150484
rect 150544 150470 151018 150498
rect 150440 147892 150492 147898
rect 150440 147834 150492 147840
rect 150452 147218 150480 147834
rect 150440 147212 150492 147218
rect 150440 147154 150492 147160
rect 150348 147076 150400 147082
rect 150348 147018 150400 147024
rect 149152 5500 149204 5506
rect 149152 5442 149204 5448
rect 149520 5228 149572 5234
rect 149520 5170 149572 5176
rect 148324 4956 148376 4962
rect 148324 4898 148376 4904
rect 147680 3868 147732 3874
rect 147680 3810 147732 3816
rect 148336 480 148364 4898
rect 149532 480 149560 5170
rect 150544 3942 150572 150470
rect 151740 147966 151768 150484
rect 151832 150470 152398 150498
rect 151728 147960 151780 147966
rect 151728 147902 151780 147908
rect 151728 13116 151780 13122
rect 151728 13058 151780 13064
rect 150532 3936 150584 3942
rect 150532 3878 150584 3884
rect 151740 3534 151768 13058
rect 151832 6186 151860 150470
rect 153120 145858 153148 150484
rect 153764 147898 153792 150484
rect 153948 150470 154514 150498
rect 153752 147892 153804 147898
rect 153752 147834 153804 147840
rect 153108 145852 153160 145858
rect 153108 145794 153160 145800
rect 153948 142154 153976 150470
rect 154856 148776 154908 148782
rect 154856 148718 154908 148724
rect 154868 147354 154896 148718
rect 154856 147348 154908 147354
rect 154856 147290 154908 147296
rect 155144 144226 155172 150484
rect 155224 148708 155276 148714
rect 155224 148650 155276 148656
rect 155132 144220 155184 144226
rect 155132 144162 155184 144168
rect 153304 142126 153976 142154
rect 153016 9240 153068 9246
rect 153016 9182 153068 9188
rect 151820 6180 151872 6186
rect 151820 6122 151872 6128
rect 151820 5092 151872 5098
rect 151820 5034 151872 5040
rect 150624 3528 150676 3534
rect 150624 3470 150676 3476
rect 151728 3528 151780 3534
rect 151728 3470 151780 3476
rect 150636 480 150664 3470
rect 151832 480 151860 5034
rect 153028 480 153056 9182
rect 153304 6254 153332 142126
rect 153292 6248 153344 6254
rect 153292 6190 153344 6196
rect 155236 4214 155264 148650
rect 155880 148034 155908 150484
rect 155972 150470 156538 150498
rect 155868 148028 155920 148034
rect 155868 147970 155920 147976
rect 155972 6322 156000 150470
rect 157260 146062 157288 150484
rect 157904 148782 157932 150484
rect 158088 150470 158562 150498
rect 158824 150470 159298 150498
rect 157892 148776 157944 148782
rect 157892 148718 157944 148724
rect 157248 146056 157300 146062
rect 157248 145998 157300 146004
rect 158088 142154 158116 150470
rect 157444 142126 158116 142154
rect 156604 9308 156656 9314
rect 156604 9250 156656 9256
rect 155960 6316 156012 6322
rect 155960 6258 156012 6264
rect 155408 5024 155460 5030
rect 155408 4966 155460 4972
rect 154212 4208 154264 4214
rect 154212 4150 154264 4156
rect 155224 4208 155276 4214
rect 155224 4150 155276 4156
rect 154224 480 154252 4150
rect 155420 480 155448 4966
rect 156616 480 156644 9250
rect 157444 6390 157472 142126
rect 158824 8974 158852 150470
rect 159928 147286 159956 150484
rect 160112 150470 160678 150498
rect 159916 147280 159968 147286
rect 159916 147222 159968 147228
rect 158812 8968 158864 8974
rect 158812 8910 158864 8916
rect 158904 8152 158956 8158
rect 158904 8094 158956 8100
rect 157432 6384 157484 6390
rect 157432 6326 157484 6332
rect 157800 5160 157852 5166
rect 157800 5102 157852 5108
rect 157812 480 157840 5102
rect 158916 480 158944 8094
rect 160112 6458 160140 150470
rect 161308 144294 161336 150484
rect 161492 150470 162058 150498
rect 162136 150470 162702 150498
rect 161296 144288 161348 144294
rect 161296 144230 161348 144236
rect 161388 18624 161440 18630
rect 161388 18566 161440 18572
rect 161296 8968 161348 8974
rect 161296 8910 161348 8916
rect 160100 6452 160152 6458
rect 160100 6394 160152 6400
rect 160100 3528 160152 3534
rect 160100 3470 160152 3476
rect 160112 480 160140 3470
rect 161308 480 161336 8910
rect 161400 3534 161428 18566
rect 161492 4758 161520 150470
rect 162136 146418 162164 150470
rect 162216 148028 162268 148034
rect 162216 147970 162268 147976
rect 161584 146390 162164 146418
rect 161584 6526 161612 146390
rect 162228 142154 162256 147970
rect 163424 145994 163452 150484
rect 163516 150470 164082 150498
rect 164252 150470 164818 150498
rect 163412 145988 163464 145994
rect 163412 145930 163464 145936
rect 163516 142154 163544 150470
rect 162136 142126 162256 142154
rect 162872 142126 163544 142154
rect 161572 6520 161624 6526
rect 161572 6462 161624 6468
rect 162136 5234 162164 142126
rect 162124 5228 162176 5234
rect 162124 5170 162176 5176
rect 162492 5228 162544 5234
rect 162492 5170 162544 5176
rect 161480 4752 161532 4758
rect 161480 4694 161532 4700
rect 161388 3528 161440 3534
rect 161388 3470 161440 3476
rect 162504 480 162532 5170
rect 162872 4622 162900 142126
rect 164252 6594 164280 150470
rect 165448 144362 165476 150484
rect 165724 150470 166106 150498
rect 165436 144356 165488 144362
rect 165436 144298 165488 144304
rect 164240 6588 164292 6594
rect 164240 6530 164292 6536
rect 164884 5296 164936 5302
rect 164884 5238 164936 5244
rect 162860 4616 162912 4622
rect 162860 4558 162912 4564
rect 163688 4208 163740 4214
rect 163688 4150 163740 4156
rect 163700 480 163728 4150
rect 164896 480 164924 5238
rect 165724 4690 165752 150470
rect 166828 148850 166856 150484
rect 166816 148844 166868 148850
rect 166816 148786 166868 148792
rect 166264 148776 166316 148782
rect 166264 148718 166316 148724
rect 166080 5364 166132 5370
rect 166080 5306 166132 5312
rect 165712 4684 165764 4690
rect 165712 4626 165764 4632
rect 166092 480 166120 5306
rect 166276 4214 166304 148718
rect 167472 146130 167500 150484
rect 167656 150470 168222 150498
rect 168484 150470 168866 150498
rect 169312 150470 169602 150498
rect 169864 150470 170246 150498
rect 167460 146124 167512 146130
rect 167460 146066 167512 146072
rect 167656 142154 167684 150470
rect 168380 144900 168432 144906
rect 168380 144842 168432 144848
rect 167012 142126 167684 142154
rect 167012 4554 167040 142126
rect 167000 4548 167052 4554
rect 167000 4490 167052 4496
rect 166264 4208 166316 4214
rect 166264 4150 166316 4156
rect 167184 4208 167236 4214
rect 167184 4150 167236 4156
rect 167196 480 167224 4150
rect 168392 4010 168420 144842
rect 168484 6662 168512 150470
rect 169312 144906 169340 150470
rect 169300 144900 169352 144906
rect 169300 144842 169352 144848
rect 169668 10328 169720 10334
rect 169668 10270 169720 10276
rect 169576 8220 169628 8226
rect 169576 8162 169628 8168
rect 168472 6656 168524 6662
rect 168472 6598 168524 6604
rect 168380 4004 168432 4010
rect 168380 3946 168432 3952
rect 168380 3528 168432 3534
rect 168380 3470 168432 3476
rect 168392 480 168420 3470
rect 169588 480 169616 8162
rect 169680 3534 169708 10270
rect 169864 4486 169892 150470
rect 170404 148096 170456 148102
rect 170404 148038 170456 148044
rect 169852 4480 169904 4486
rect 169852 4422 169904 4428
rect 170416 4214 170444 148038
rect 170968 147966 170996 150484
rect 171152 150470 171626 150498
rect 171704 150470 172362 150498
rect 172624 150470 173006 150498
rect 173084 150470 173742 150498
rect 174004 150470 174386 150498
rect 170956 147960 171008 147966
rect 170956 147902 171008 147908
rect 170772 6180 170824 6186
rect 170772 6122 170824 6128
rect 170404 4208 170456 4214
rect 170404 4150 170456 4156
rect 169668 3528 169720 3534
rect 169668 3470 169720 3476
rect 170784 480 170812 6122
rect 171152 4078 171180 150470
rect 171704 142154 171732 150470
rect 171244 142126 171732 142154
rect 171244 4418 171272 142126
rect 172624 6730 172652 150470
rect 173084 142154 173112 150470
rect 173164 148844 173216 148850
rect 173164 148786 173216 148792
rect 172716 142126 173112 142154
rect 172612 6724 172664 6730
rect 172612 6666 172664 6672
rect 171232 4412 171284 4418
rect 171232 4354 171284 4360
rect 171968 4208 172020 4214
rect 171968 4150 172020 4156
rect 171140 4072 171192 4078
rect 171140 4014 171192 4020
rect 171980 480 172008 4150
rect 172716 3398 172744 142126
rect 173176 4214 173204 148786
rect 173256 6248 173308 6254
rect 173256 6190 173308 6196
rect 173164 4208 173216 4214
rect 173164 4150 173216 4156
rect 172704 3392 172756 3398
rect 172704 3334 172756 3340
rect 173268 3176 173296 6190
rect 174004 4350 174032 150470
rect 175016 147422 175044 150484
rect 175292 150470 175766 150498
rect 176120 150470 176410 150498
rect 175004 147416 175056 147422
rect 175004 147358 175056 147364
rect 174268 8288 174320 8294
rect 174268 8230 174320 8236
rect 173992 4344 174044 4350
rect 173992 4286 174044 4292
rect 173176 3148 173296 3176
rect 173176 480 173204 3148
rect 174280 480 174308 8230
rect 175292 4146 175320 150470
rect 176120 142154 176148 150470
rect 177132 148918 177160 150484
rect 177224 150470 177790 150498
rect 177120 148912 177172 148918
rect 177120 148854 177172 148860
rect 177224 142154 177252 150470
rect 177304 148912 177356 148918
rect 177304 148854 177356 148860
rect 177316 147558 177344 148854
rect 177304 147552 177356 147558
rect 177304 147494 177356 147500
rect 178512 147490 178540 150484
rect 178880 150470 179170 150498
rect 179616 150470 179906 150498
rect 180168 150470 180550 150498
rect 178500 147484 178552 147490
rect 178500 147426 178552 147432
rect 178880 142154 178908 150470
rect 179512 146328 179564 146334
rect 179512 146270 179564 146276
rect 175384 142126 176148 142154
rect 176856 142126 177252 142154
rect 178144 142126 178908 142154
rect 175384 4282 175412 142126
rect 175464 4752 175516 4758
rect 175464 4694 175516 4700
rect 175372 4276 175424 4282
rect 175372 4218 175424 4224
rect 175280 4140 175332 4146
rect 175280 4082 175332 4088
rect 175476 480 175504 4694
rect 176660 3528 176712 3534
rect 176660 3470 176712 3476
rect 176672 480 176700 3470
rect 176856 3330 176884 142126
rect 177948 14476 178000 14482
rect 177948 14418 178000 14424
rect 177856 6316 177908 6322
rect 177856 6258 177908 6264
rect 176844 3324 176896 3330
rect 176844 3266 176896 3272
rect 177868 480 177896 6258
rect 177960 3534 177988 14418
rect 178144 9042 178172 142126
rect 178132 9036 178184 9042
rect 178132 8978 178184 8984
rect 179524 6798 179552 146270
rect 179512 6792 179564 6798
rect 179512 6734 179564 6740
rect 179052 6384 179104 6390
rect 179052 6326 179104 6332
rect 177948 3528 178000 3534
rect 177948 3470 178000 3476
rect 179064 480 179092 6326
rect 179616 3262 179644 150470
rect 180168 146334 180196 150470
rect 181272 148918 181300 150484
rect 181364 150470 181930 150498
rect 182284 150470 182574 150498
rect 181260 148912 181312 148918
rect 181260 148854 181312 148860
rect 180156 146328 180208 146334
rect 180156 146270 180208 146276
rect 181364 142154 181392 150470
rect 180996 142126 181392 142154
rect 180708 17264 180760 17270
rect 180708 17206 180760 17212
rect 180720 3534 180748 17206
rect 180248 3528 180300 3534
rect 180248 3470 180300 3476
rect 180708 3528 180760 3534
rect 180708 3470 180760 3476
rect 179604 3256 179656 3262
rect 179604 3198 179656 3204
rect 180260 480 180288 3470
rect 180996 3194 181024 142126
rect 182284 6118 182312 150470
rect 183296 148986 183324 150484
rect 183756 150470 183954 150498
rect 184400 150470 184690 150498
rect 183284 148980 183336 148986
rect 183284 148922 183336 148928
rect 183652 146328 183704 146334
rect 183652 146270 183704 146276
rect 182272 6112 182324 6118
rect 182272 6054 182324 6060
rect 183664 6050 183692 146270
rect 183756 16574 183784 150470
rect 184204 148912 184256 148918
rect 184204 148854 184256 148860
rect 183756 16546 183876 16574
rect 183744 6452 183796 6458
rect 183744 6394 183796 6400
rect 183652 6044 183704 6050
rect 183652 5986 183704 5992
rect 182548 4208 182600 4214
rect 182548 4150 182600 4156
rect 181444 3460 181496 3466
rect 181444 3402 181496 3408
rect 180984 3188 181036 3194
rect 180984 3130 181036 3136
rect 181456 480 181484 3402
rect 182560 480 182588 4150
rect 183756 480 183784 6394
rect 183848 3126 183876 16546
rect 184216 4214 184244 148854
rect 184400 146334 184428 150470
rect 185320 147694 185348 150484
rect 186056 149054 186084 150484
rect 186424 150470 186714 150498
rect 186044 149048 186096 149054
rect 186044 148990 186096 148996
rect 185308 147688 185360 147694
rect 185308 147630 185360 147636
rect 184388 146328 184440 146334
rect 184388 146270 184440 146276
rect 186424 5982 186452 150470
rect 187436 148306 187464 150484
rect 187712 150470 188094 150498
rect 188356 150470 188830 150498
rect 189092 150470 189474 150498
rect 187608 148980 187660 148986
rect 187608 148922 187660 148928
rect 187424 148300 187476 148306
rect 187424 148242 187476 148248
rect 187620 6914 187648 148922
rect 187344 6886 187648 6914
rect 186412 5976 186464 5982
rect 186412 5918 186464 5924
rect 186136 5432 186188 5438
rect 186136 5374 186188 5380
rect 184204 4208 184256 4214
rect 184204 4150 184256 4156
rect 184940 3528 184992 3534
rect 184940 3470 184992 3476
rect 183836 3120 183888 3126
rect 183836 3062 183888 3068
rect 184952 480 184980 3470
rect 186148 480 186176 5374
rect 187344 480 187372 6886
rect 187712 3058 187740 150470
rect 188356 142154 188384 150470
rect 189092 147778 189120 150470
rect 190196 148238 190224 150484
rect 190564 150470 190854 150498
rect 190184 148232 190236 148238
rect 190184 148174 190236 148180
rect 189000 147750 189120 147778
rect 189000 146878 189028 147750
rect 188988 146872 189040 146878
rect 188988 146814 189040 146820
rect 187804 142126 188384 142154
rect 187804 5914 187832 142126
rect 187792 5908 187844 5914
rect 187792 5850 187844 5856
rect 190564 5846 190592 150470
rect 191484 148170 191512 150484
rect 191852 150470 192234 150498
rect 192312 150470 192878 150498
rect 191748 149048 191800 149054
rect 191748 148990 191800 148996
rect 191472 148164 191524 148170
rect 191472 148106 191524 148112
rect 191104 147688 191156 147694
rect 191104 147630 191156 147636
rect 191116 141438 191144 147630
rect 191104 141432 191156 141438
rect 191104 141374 191156 141380
rect 190552 5840 190604 5846
rect 190552 5782 190604 5788
rect 189724 5500 189776 5506
rect 189724 5442 189776 5448
rect 188528 3596 188580 3602
rect 188528 3538 188580 3544
rect 187700 3052 187752 3058
rect 187700 2994 187752 3000
rect 188540 480 188568 3538
rect 189736 480 189764 5442
rect 191760 3058 191788 148990
rect 190828 3052 190880 3058
rect 190828 2994 190880 3000
rect 191748 3052 191800 3058
rect 191748 2994 191800 3000
rect 190840 480 190868 2994
rect 191852 2990 191880 150470
rect 192312 142154 192340 150470
rect 193600 147694 193628 150484
rect 193876 150470 194258 150498
rect 194612 150470 194994 150498
rect 193588 147688 193640 147694
rect 193588 147630 193640 147636
rect 193876 142154 193904 150470
rect 191944 142126 192340 142154
rect 193416 142126 193904 142154
rect 191944 5778 191972 142126
rect 191932 5772 191984 5778
rect 191932 5714 191984 5720
rect 193220 4208 193272 4214
rect 193220 4150 193272 4156
rect 192024 3732 192076 3738
rect 192024 3674 192076 3680
rect 191840 2984 191892 2990
rect 191840 2926 191892 2932
rect 192036 480 192064 3674
rect 193232 480 193260 4150
rect 193416 2922 193444 142126
rect 194612 5710 194640 150470
rect 195244 148300 195296 148306
rect 195244 148242 195296 148248
rect 194600 5704 194652 5710
rect 194600 5646 194652 5652
rect 194416 4276 194468 4282
rect 194416 4218 194468 4224
rect 193404 2916 193456 2922
rect 193404 2858 193456 2864
rect 194428 480 194456 4218
rect 195256 4214 195284 148242
rect 195624 146198 195652 150484
rect 196176 150470 196374 150498
rect 196728 150470 197018 150498
rect 197464 150470 197754 150498
rect 196072 146328 196124 146334
rect 196072 146270 196124 146276
rect 195612 146192 195664 146198
rect 195612 146134 195664 146140
rect 196084 7614 196112 146270
rect 196072 7608 196124 7614
rect 196072 7550 196124 7556
rect 195244 4208 195296 4214
rect 195244 4150 195296 4156
rect 195612 3664 195664 3670
rect 195612 3606 195664 3612
rect 195624 480 195652 3606
rect 196176 2854 196204 150470
rect 196624 148232 196676 148238
rect 196624 148174 196676 148180
rect 196636 4758 196664 148174
rect 196728 146334 196756 150470
rect 196716 146328 196768 146334
rect 196716 146270 196768 146276
rect 197464 7682 197492 150470
rect 198384 148374 198412 150484
rect 199028 148510 199056 150484
rect 199120 150470 199778 150498
rect 199016 148504 199068 148510
rect 199016 148446 199068 148452
rect 198372 148368 198424 148374
rect 198372 148310 198424 148316
rect 198004 148164 198056 148170
rect 198004 148106 198056 148112
rect 197452 7676 197504 7682
rect 197452 7618 197504 7624
rect 196808 7608 196860 7614
rect 196808 7550 196860 7556
rect 196624 4752 196676 4758
rect 196624 4694 196676 4700
rect 196164 2848 196216 2854
rect 196164 2790 196216 2796
rect 196820 480 196848 7550
rect 198016 4282 198044 148106
rect 199120 142154 199148 150470
rect 200408 148442 200436 150484
rect 200592 150470 201158 150498
rect 201604 150470 201802 150498
rect 202248 150470 202538 150498
rect 200396 148436 200448 148442
rect 200396 148378 200448 148384
rect 200592 142154 200620 150470
rect 200764 147756 200816 147762
rect 200764 147698 200816 147704
rect 198844 142126 199148 142154
rect 200224 142126 200620 142154
rect 198844 7750 198872 142126
rect 200224 11762 200252 142126
rect 200212 11756 200264 11762
rect 200212 11698 200264 11704
rect 200776 8022 200804 147698
rect 201500 146328 201552 146334
rect 201500 146270 201552 146276
rect 200764 8016 200816 8022
rect 200764 7958 200816 7964
rect 201512 7886 201540 146270
rect 201500 7880 201552 7886
rect 201500 7822 201552 7828
rect 201604 7818 201632 150470
rect 202144 147688 202196 147694
rect 202144 147630 202196 147636
rect 202156 15910 202184 147630
rect 202248 146334 202276 150470
rect 203168 148646 203196 150484
rect 203156 148640 203208 148646
rect 203156 148582 203208 148588
rect 203904 147694 203932 150484
rect 204548 147762 204576 150484
rect 204640 150470 205298 150498
rect 205652 150470 205942 150498
rect 206112 150470 206678 150498
rect 204536 147756 204588 147762
rect 204536 147698 204588 147704
rect 203892 147688 203944 147694
rect 203892 147630 203944 147636
rect 202236 146328 202288 146334
rect 202236 146270 202288 146276
rect 204640 142154 204668 150470
rect 205548 148368 205600 148374
rect 205548 148310 205600 148316
rect 204364 142126 204668 142154
rect 202144 15904 202196 15910
rect 202144 15846 202196 15852
rect 204364 7954 204392 142126
rect 204352 7948 204404 7954
rect 204352 7890 204404 7896
rect 201592 7812 201644 7818
rect 201592 7754 201644 7760
rect 198832 7744 198884 7750
rect 198832 7686 198884 7692
rect 203892 4752 203944 4758
rect 203892 4694 203944 4700
rect 200304 4684 200356 4690
rect 200304 4626 200356 4632
rect 198004 4276 198056 4282
rect 198004 4218 198056 4224
rect 199108 3868 199160 3874
rect 199108 3810 199160 3816
rect 197912 3800 197964 3806
rect 197912 3742 197964 3748
rect 197924 480 197952 3742
rect 199120 480 199148 3810
rect 200316 480 200344 4626
rect 201500 4004 201552 4010
rect 201500 3946 201552 3952
rect 201512 480 201540 3946
rect 202696 3936 202748 3942
rect 202696 3878 202748 3884
rect 202708 480 202736 3878
rect 203904 480 203932 4694
rect 205560 3398 205588 148310
rect 205652 4826 205680 150470
rect 206112 142154 206140 150470
rect 207308 148578 207336 150484
rect 207400 150470 207966 150498
rect 208504 150470 208702 150498
rect 209056 150470 209346 150498
rect 209884 150470 210082 150498
rect 207296 148572 207348 148578
rect 207296 148514 207348 148520
rect 207400 142154 207428 150470
rect 208400 147824 208452 147830
rect 208400 147766 208452 147772
rect 205744 142126 206140 142154
rect 207124 142126 207428 142154
rect 205744 9178 205772 142126
rect 205732 9172 205784 9178
rect 205732 9114 205784 9120
rect 207124 4894 207152 142126
rect 208412 8090 208440 147766
rect 208504 9110 208532 150470
rect 209056 147830 209084 150470
rect 209044 147824 209096 147830
rect 209044 147766 209096 147772
rect 209044 147688 209096 147694
rect 209044 147630 209096 147636
rect 209056 13122 209084 147630
rect 209044 13116 209096 13122
rect 209044 13058 209096 13064
rect 208492 9104 208544 9110
rect 208492 9046 208544 9052
rect 208400 8084 208452 8090
rect 208400 8026 208452 8032
rect 209884 4962 209912 150470
rect 210712 148034 210740 150484
rect 210700 148028 210752 148034
rect 210700 147970 210752 147976
rect 211448 147694 211476 150484
rect 211816 150470 212106 150498
rect 212644 150470 212842 150498
rect 211436 147688 211488 147694
rect 211436 147630 211488 147636
rect 211816 142154 211844 150470
rect 211264 142126 211844 142154
rect 211264 5098 211292 142126
rect 212644 9246 212672 150470
rect 213472 148714 213500 150484
rect 213932 150470 214222 150498
rect 214576 150470 214866 150498
rect 215312 150470 215510 150498
rect 215772 150470 216246 150498
rect 216784 150470 216890 150498
rect 217336 150470 217626 150498
rect 218164 150470 218270 150498
rect 213460 148708 213512 148714
rect 213460 148650 213512 148656
rect 213828 148436 213880 148442
rect 213828 148378 213880 148384
rect 212632 9240 212684 9246
rect 212632 9182 212684 9188
rect 211252 5092 211304 5098
rect 211252 5034 211304 5040
rect 209872 4956 209924 4962
rect 209872 4898 209924 4904
rect 207112 4888 207164 4894
rect 207112 4830 207164 4836
rect 210976 4888 211028 4894
rect 210976 4830 211028 4836
rect 205640 4820 205692 4826
rect 205640 4762 205692 4768
rect 207388 4820 207440 4826
rect 207388 4762 207440 4768
rect 206192 4072 206244 4078
rect 206192 4014 206244 4020
rect 205088 3392 205140 3398
rect 205088 3334 205140 3340
rect 205548 3392 205600 3398
rect 205548 3334 205600 3340
rect 205100 480 205128 3334
rect 206204 480 206232 4014
rect 207400 480 207428 4762
rect 208584 4140 208636 4146
rect 208584 4082 208636 4088
rect 208596 480 208624 4082
rect 209780 3256 209832 3262
rect 209780 3198 209832 3204
rect 209792 480 209820 3198
rect 210988 480 211016 4830
rect 213840 3398 213868 148378
rect 213932 5030 213960 150470
rect 214576 142154 214604 150470
rect 214024 142126 214604 142154
rect 214024 9314 214052 142126
rect 215208 15904 215260 15910
rect 215208 15846 215260 15852
rect 214012 9308 214064 9314
rect 214012 9250 214064 9256
rect 213920 5024 213972 5030
rect 213920 4966 213972 4972
rect 215220 3398 215248 15846
rect 215312 5166 215340 150470
rect 215772 142154 215800 150470
rect 216680 146328 216732 146334
rect 216680 146270 216732 146276
rect 215404 142126 215800 142154
rect 215404 8158 215432 142126
rect 216692 8974 216720 146270
rect 216784 18630 216812 150470
rect 217336 146334 217364 150470
rect 217324 146328 217376 146334
rect 217324 146270 217376 146276
rect 216772 18624 216824 18630
rect 216772 18566 216824 18572
rect 216680 8968 216732 8974
rect 216680 8910 216732 8916
rect 215392 8152 215444 8158
rect 215392 8094 215444 8100
rect 218164 5234 218192 150470
rect 218992 148782 219020 150484
rect 219544 150470 219650 150498
rect 220096 150470 220386 150498
rect 218980 148776 219032 148782
rect 218980 148718 219032 148724
rect 219440 147824 219492 147830
rect 219440 147766 219492 147772
rect 219452 5370 219480 147766
rect 219440 5364 219492 5370
rect 219440 5306 219492 5312
rect 219544 5302 219572 150470
rect 220096 147830 220124 150470
rect 221016 148102 221044 150484
rect 221004 148096 221056 148102
rect 221004 148038 221056 148044
rect 220084 147824 220136 147830
rect 220084 147766 220136 147772
rect 221752 147694 221780 150484
rect 222304 150470 222410 150498
rect 222856 150470 223146 150498
rect 220084 147688 220136 147694
rect 220084 147630 220136 147636
rect 221740 147688 221792 147694
rect 221740 147630 221792 147636
rect 220096 10334 220124 147630
rect 222200 146328 222252 146334
rect 222200 146270 222252 146276
rect 220084 10328 220136 10334
rect 220084 10270 220136 10276
rect 222212 6186 222240 146270
rect 222304 8226 222332 150470
rect 222856 146334 222884 150470
rect 223776 148850 223804 150484
rect 224144 150470 224434 150498
rect 223764 148844 223816 148850
rect 223764 148786 223816 148792
rect 223488 148572 223540 148578
rect 223488 148514 223540 148520
rect 222844 146328 222896 146334
rect 222844 146270 222896 146276
rect 222292 8220 222344 8226
rect 222292 8162 222344 8168
rect 222200 6180 222252 6186
rect 222200 6122 222252 6128
rect 219532 5296 219584 5302
rect 219532 5238 219584 5244
rect 218152 5228 218204 5234
rect 218152 5170 218204 5176
rect 215300 5160 215352 5166
rect 215300 5102 215352 5108
rect 218060 5024 218112 5030
rect 218060 4966 218112 4972
rect 213368 3392 213420 3398
rect 213368 3334 213420 3340
rect 213828 3392 213880 3398
rect 213828 3334 213880 3340
rect 214472 3392 214524 3398
rect 214472 3334 214524 3340
rect 215208 3392 215260 3398
rect 215208 3334 215260 3340
rect 212172 3188 212224 3194
rect 212172 3130 212224 3136
rect 212184 480 212212 3130
rect 213380 480 213408 3334
rect 214484 480 214512 3334
rect 216864 3188 216916 3194
rect 216864 3130 216916 3136
rect 215668 3120 215720 3126
rect 215668 3062 215720 3068
rect 215680 480 215708 3062
rect 216876 480 216904 3130
rect 218072 480 218100 4966
rect 221556 4956 221608 4962
rect 221556 4898 221608 4904
rect 219256 3256 219308 3262
rect 219256 3198 219308 3204
rect 219268 480 219296 3198
rect 220452 2984 220504 2990
rect 220452 2926 220504 2932
rect 220464 480 220492 2926
rect 221568 480 221596 4898
rect 223500 3058 223528 148514
rect 224144 142154 224172 150470
rect 224868 148504 224920 148510
rect 224868 148446 224920 148452
rect 224224 147688 224276 147694
rect 224224 147630 224276 147636
rect 223684 142126 224172 142154
rect 223684 6254 223712 142126
rect 224236 8294 224264 147630
rect 224224 8288 224276 8294
rect 224224 8230 224276 8236
rect 223672 6248 223724 6254
rect 223672 6190 223724 6196
rect 224880 3058 224908 148446
rect 225156 147694 225184 150484
rect 225800 148238 225828 150484
rect 226444 150470 226550 150498
rect 226904 150470 227194 150498
rect 227732 150470 227930 150498
rect 228100 150470 228574 150498
rect 225788 148232 225840 148238
rect 225788 148174 225840 148180
rect 225144 147688 225196 147694
rect 225144 147630 225196 147636
rect 226340 146328 226392 146334
rect 226340 146270 226392 146276
rect 226352 6322 226380 146270
rect 226444 14482 226472 150470
rect 226904 146334 226932 150470
rect 227628 148640 227680 148646
rect 227628 148582 227680 148588
rect 226892 146328 226944 146334
rect 226892 146270 226944 146276
rect 226432 14476 226484 14482
rect 226432 14418 226484 14424
rect 226340 6316 226392 6322
rect 226340 6258 226392 6264
rect 226524 3664 226576 3670
rect 226524 3606 226576 3612
rect 226536 3534 226564 3606
rect 226524 3528 226576 3534
rect 226524 3470 226576 3476
rect 222752 3052 222804 3058
rect 222752 2994 222804 3000
rect 223488 3052 223540 3058
rect 223488 2994 223540 3000
rect 223948 3052 224000 3058
rect 223948 2994 224000 3000
rect 224868 3052 224920 3058
rect 224868 2994 224920 3000
rect 226340 3052 226392 3058
rect 226340 2994 226392 3000
rect 222764 480 222792 2994
rect 223960 480 223988 2994
rect 225144 2916 225196 2922
rect 225144 2858 225196 2864
rect 225156 480 225184 2858
rect 226352 480 226380 2994
rect 227640 2774 227668 148582
rect 227732 6390 227760 150470
rect 228100 142154 228128 150470
rect 228364 148232 228416 148238
rect 228364 148174 228416 148180
rect 227824 142126 228128 142154
rect 227824 17270 227852 142126
rect 227812 17264 227864 17270
rect 227812 17206 227864 17212
rect 227720 6384 227772 6390
rect 227720 6326 227772 6332
rect 228376 4690 228404 148174
rect 228364 4684 228416 4690
rect 228364 4626 228416 4632
rect 229296 3466 229324 150484
rect 229940 148918 229968 150484
rect 230584 150470 230690 150498
rect 230952 150470 231334 150498
rect 229928 148912 229980 148918
rect 229928 148854 229980 148860
rect 230584 6458 230612 150470
rect 230952 142154 230980 150470
rect 231768 148708 231820 148714
rect 231768 148650 231820 148656
rect 230676 142126 230980 142154
rect 230572 6452 230624 6458
rect 230572 6394 230624 6400
rect 229836 3868 229888 3874
rect 229888 3828 229968 3856
rect 229836 3810 229888 3816
rect 229940 3738 229968 3828
rect 229928 3732 229980 3738
rect 229928 3674 229980 3680
rect 229836 3664 229888 3670
rect 229836 3606 229888 3612
rect 229284 3460 229336 3466
rect 229284 3402 229336 3408
rect 228732 2848 228784 2854
rect 228732 2790 228784 2796
rect 227548 2746 227668 2774
rect 227548 480 227576 2746
rect 228744 480 228772 2790
rect 229848 480 229876 3606
rect 230676 3466 230704 142126
rect 231780 3874 231808 148650
rect 231964 5438 231992 150484
rect 232700 148986 232728 150484
rect 232688 148980 232740 148986
rect 232688 148922 232740 148928
rect 232504 147688 232556 147694
rect 232504 147630 232556 147636
rect 232516 5506 232544 147630
rect 232504 5500 232556 5506
rect 232504 5442 232556 5448
rect 231952 5432 232004 5438
rect 231952 5374 232004 5380
rect 231032 3868 231084 3874
rect 231032 3810 231084 3816
rect 231768 3868 231820 3874
rect 231768 3810 231820 3816
rect 230664 3460 230716 3466
rect 230664 3402 230716 3408
rect 231044 480 231072 3810
rect 233344 3534 233372 150484
rect 234080 147694 234108 150484
rect 234724 149054 234752 150484
rect 235000 150470 235474 150498
rect 234712 149048 234764 149054
rect 234712 148990 234764 148996
rect 234528 148776 234580 148782
rect 234528 148718 234580 148724
rect 234068 147688 234120 147694
rect 234068 147630 234120 147636
rect 234540 3534 234568 148718
rect 235000 142154 235028 150470
rect 235908 148980 235960 148986
rect 235908 148922 235960 148928
rect 234724 142126 235028 142154
rect 234724 3602 234752 142126
rect 234712 3596 234764 3602
rect 234712 3538 234764 3544
rect 235816 3596 235868 3602
rect 235816 3538 235868 3544
rect 233332 3528 233384 3534
rect 233332 3470 233384 3476
rect 233424 3528 233476 3534
rect 233424 3470 233476 3476
rect 234528 3528 234580 3534
rect 234528 3470 234580 3476
rect 234620 3528 234672 3534
rect 234620 3470 234672 3476
rect 232228 3460 232280 3466
rect 232228 3402 232280 3408
rect 232240 480 232268 3402
rect 233436 480 233464 3470
rect 234632 480 234660 3470
rect 235828 480 235856 3538
rect 235920 3534 235948 148922
rect 236104 148306 236132 150484
rect 236092 148300 236144 148306
rect 236092 148242 236144 148248
rect 236840 148170 236868 150484
rect 237392 150470 237498 150498
rect 237760 150470 238234 150498
rect 238772 150470 238878 150498
rect 239140 150470 239614 150498
rect 237288 148844 237340 148850
rect 237288 148786 237340 148792
rect 236828 148164 236880 148170
rect 236828 148106 236880 148112
rect 237300 6914 237328 148786
rect 237024 6886 237328 6914
rect 235908 3528 235960 3534
rect 235908 3470 235960 3476
rect 237024 480 237052 6886
rect 237392 3874 237420 150470
rect 237760 142154 237788 150470
rect 238668 148912 238720 148918
rect 238668 148854 238720 148860
rect 237484 142126 237788 142154
rect 237484 7614 237512 142126
rect 237472 7608 237524 7614
rect 237472 7550 237524 7556
rect 237380 3868 237432 3874
rect 237380 3810 237432 3816
rect 238680 3670 238708 148854
rect 238772 3806 238800 150470
rect 239140 142154 239168 150470
rect 240244 148238 240272 150484
rect 240428 150470 240902 150498
rect 241532 150470 241638 150498
rect 241808 150470 242282 150498
rect 240232 148232 240284 148238
rect 240232 148174 240284 148180
rect 240428 142154 240456 150470
rect 241428 149048 241480 149054
rect 241428 148990 241480 148996
rect 240784 148096 240836 148102
rect 240784 148038 240836 148044
rect 238864 142126 239168 142154
rect 240244 142126 240456 142154
rect 238760 3800 238812 3806
rect 238760 3742 238812 3748
rect 238864 3738 238892 142126
rect 240244 3874 240272 142126
rect 240796 5030 240824 148038
rect 240784 5024 240836 5030
rect 240784 4966 240836 4972
rect 240232 3868 240284 3874
rect 240232 3810 240284 3816
rect 238852 3732 238904 3738
rect 238852 3674 238904 3680
rect 239312 3732 239364 3738
rect 239312 3674 239364 3680
rect 238116 3664 238168 3670
rect 238116 3606 238168 3612
rect 238668 3664 238720 3670
rect 238668 3606 238720 3612
rect 238128 480 238156 3606
rect 239324 480 239352 3674
rect 241440 3466 241468 148990
rect 241532 4010 241560 150470
rect 241808 142154 241836 150470
rect 243004 148374 243032 150484
rect 243280 150470 243662 150498
rect 242992 148368 243044 148374
rect 242992 148310 243044 148316
rect 242808 148300 242860 148306
rect 242808 148242 242860 148248
rect 241624 142126 241836 142154
rect 241624 4758 241652 142126
rect 241612 4752 241664 4758
rect 241612 4694 241664 4700
rect 241520 4004 241572 4010
rect 241520 3946 241572 3952
rect 242820 3466 242848 148242
rect 243280 142154 243308 150470
rect 244188 148164 244240 148170
rect 244188 148106 244240 148112
rect 243004 142126 243308 142154
rect 243004 4078 243032 142126
rect 242992 4072 243044 4078
rect 242992 4014 243044 4020
rect 244200 3466 244228 148106
rect 244280 145716 244332 145722
rect 244280 145658 244332 145664
rect 244292 4146 244320 145658
rect 244384 4826 244412 150484
rect 244752 150470 245042 150498
rect 245672 150470 245778 150498
rect 245856 150470 246422 150498
rect 247158 150470 247264 150498
rect 244752 145722 244780 150470
rect 244924 148368 244976 148374
rect 244924 148310 244976 148316
rect 244740 145716 244792 145722
rect 244740 145658 244792 145664
rect 244372 4820 244424 4826
rect 244372 4762 244424 4768
rect 244280 4140 244332 4146
rect 244280 4082 244332 4088
rect 240508 3460 240560 3466
rect 240508 3402 240560 3408
rect 241428 3460 241480 3466
rect 241428 3402 241480 3408
rect 241704 3460 241756 3466
rect 241704 3402 241756 3408
rect 242808 3460 242860 3466
rect 242808 3402 242860 3408
rect 242900 3460 242952 3466
rect 242900 3402 242952 3408
rect 244188 3460 244240 3466
rect 244188 3402 244240 3408
rect 240520 480 240548 3402
rect 241716 480 241744 3402
rect 242912 480 242940 3402
rect 244936 3398 244964 148310
rect 245672 142186 245700 150470
rect 245856 146418 245884 150470
rect 246948 148232 247000 148238
rect 246948 148174 247000 148180
rect 245764 146390 245884 146418
rect 245660 142180 245712 142186
rect 245660 142122 245712 142128
rect 245764 4894 245792 146390
rect 245844 142180 245896 142186
rect 245844 142122 245896 142128
rect 245752 4888 245804 4894
rect 245752 4830 245804 4836
rect 245200 3800 245252 3806
rect 245200 3742 245252 3748
rect 244096 3392 244148 3398
rect 244096 3334 244148 3340
rect 244924 3392 244976 3398
rect 244924 3334 244976 3340
rect 244108 480 244136 3334
rect 245212 480 245240 3742
rect 245856 3670 245884 142122
rect 245844 3664 245896 3670
rect 245844 3606 245896 3612
rect 246960 3466 246988 148174
rect 247236 3942 247264 150470
rect 247788 148442 247816 150484
rect 248446 150470 248552 150498
rect 247776 148436 247828 148442
rect 247776 148378 247828 148384
rect 248524 15910 248552 150470
rect 248616 150470 249182 150498
rect 249826 150470 249932 150498
rect 248512 15904 248564 15910
rect 248512 15846 248564 15852
rect 247224 3936 247276 3942
rect 247224 3878 247276 3884
rect 247592 3664 247644 3670
rect 247592 3606 247644 3612
rect 246396 3460 246448 3466
rect 246396 3402 246448 3408
rect 246948 3460 247000 3466
rect 246948 3402 247000 3408
rect 246408 480 246436 3402
rect 247604 480 247632 3606
rect 248616 3126 248644 150470
rect 249708 148436 249760 148442
rect 249708 148378 249760 148384
rect 249720 3466 249748 148378
rect 248788 3460 248840 3466
rect 248788 3402 248840 3408
rect 249708 3460 249760 3466
rect 249708 3402 249760 3408
rect 248604 3120 248656 3126
rect 248604 3062 248656 3068
rect 248800 480 248828 3402
rect 249904 3194 249932 150470
rect 250548 148102 250576 150484
rect 251206 150470 251312 150498
rect 250536 148096 250588 148102
rect 250536 148038 250588 148044
rect 251088 148028 251140 148034
rect 251088 147970 251140 147976
rect 250444 147756 250496 147762
rect 250444 147698 250496 147704
rect 250456 3738 250484 147698
rect 250444 3732 250496 3738
rect 250444 3674 250496 3680
rect 251100 3466 251128 147970
rect 249984 3460 250036 3466
rect 249984 3402 250036 3408
rect 251088 3460 251140 3466
rect 251088 3402 251140 3408
rect 251180 3460 251232 3466
rect 251180 3402 251232 3408
rect 249892 3188 249944 3194
rect 249892 3130 249944 3136
rect 249996 480 250024 3402
rect 251192 480 251220 3402
rect 251284 3262 251312 150470
rect 251468 150470 251942 150498
rect 252586 150470 252692 150498
rect 251272 3256 251324 3262
rect 251272 3198 251324 3204
rect 251468 3058 251496 150470
rect 252468 148096 252520 148102
rect 252468 148038 252520 148044
rect 252376 3732 252428 3738
rect 252376 3674 252428 3680
rect 251456 3052 251508 3058
rect 251456 2994 251508 3000
rect 252388 480 252416 3674
rect 252480 3466 252508 148038
rect 252664 4962 252692 150470
rect 253308 148578 253336 150484
rect 253296 148572 253348 148578
rect 253296 148514 253348 148520
rect 253848 148572 253900 148578
rect 253848 148514 253900 148520
rect 253204 147824 253256 147830
rect 253204 147766 253256 147772
rect 252652 4956 252704 4962
rect 252652 4898 252704 4904
rect 253216 3806 253244 147766
rect 253204 3800 253256 3806
rect 253204 3742 253256 3748
rect 252468 3460 252520 3466
rect 252468 3402 252520 3408
rect 253492 598 253704 626
rect 253492 480 253520 598
rect 253676 490 253704 598
rect 253860 490 253888 148514
rect 253952 148510 253980 150484
rect 254136 150470 254702 150498
rect 255346 150470 255452 150498
rect 253940 148504 253992 148510
rect 253940 148446 253992 148452
rect 254136 2922 254164 150470
rect 254676 3392 254728 3398
rect 254676 3334 254728 3340
rect 254124 2916 254176 2922
rect 254124 2858 254176 2864
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 253676 462 253888 490
rect 254688 480 254716 3334
rect 255424 2990 255452 150470
rect 256068 148646 256096 150484
rect 256056 148640 256108 148646
rect 256056 148582 256108 148588
rect 256608 148504 256660 148510
rect 256608 148446 256660 148452
rect 255964 147960 256016 147966
rect 255964 147902 256016 147908
rect 255872 3460 255924 3466
rect 255872 3402 255924 3408
rect 255412 2984 255464 2990
rect 255412 2926 255464 2932
rect 255884 480 255912 3402
rect 255976 3398 256004 147902
rect 256620 3466 256648 148446
rect 256712 142186 256740 150484
rect 256804 150470 257370 150498
rect 256700 142180 256752 142186
rect 256700 142122 256752 142128
rect 256608 3460 256660 3466
rect 256608 3402 256660 3408
rect 255964 3392 256016 3398
rect 255964 3334 256016 3340
rect 256804 3330 256832 150470
rect 258092 148714 258120 150484
rect 258184 150470 258750 150498
rect 258080 148708 258132 148714
rect 258080 148650 258132 148656
rect 257988 147892 258040 147898
rect 257988 147834 258040 147840
rect 256884 142180 256936 142186
rect 256884 142122 256936 142128
rect 256792 3324 256844 3330
rect 256792 3266 256844 3272
rect 256896 2854 256924 142122
rect 258000 3466 258028 147834
rect 258184 3534 258212 150470
rect 259472 148782 259500 150484
rect 260116 148986 260144 150484
rect 260866 150470 260972 150498
rect 260104 148980 260156 148986
rect 260104 148922 260156 148928
rect 260748 148980 260800 148986
rect 260748 148922 260800 148928
rect 259460 148776 259512 148782
rect 259460 148718 259512 148724
rect 259368 148708 259420 148714
rect 259368 148650 259420 148656
rect 259380 3534 259408 148650
rect 260656 148640 260708 148646
rect 260656 148582 260708 148588
rect 258172 3528 258224 3534
rect 258172 3470 258224 3476
rect 258264 3528 258316 3534
rect 258264 3470 258316 3476
rect 259368 3528 259420 3534
rect 259368 3470 259420 3476
rect 259460 3528 259512 3534
rect 259460 3470 259512 3476
rect 257068 3460 257120 3466
rect 257068 3402 257120 3408
rect 257988 3460 258040 3466
rect 257988 3402 258040 3408
rect 256884 2848 256936 2854
rect 256884 2790 256936 2796
rect 257080 480 257108 3402
rect 258276 480 258304 3470
rect 259472 480 259500 3470
rect 260668 480 260696 148582
rect 260760 3534 260788 148922
rect 260944 3602 260972 150470
rect 261496 148850 261524 150484
rect 262232 148918 262260 150484
rect 262600 150470 262890 150498
rect 262220 148912 262272 148918
rect 262220 148854 262272 148860
rect 261484 148844 261536 148850
rect 261484 148786 261536 148792
rect 262600 147762 262628 150470
rect 263612 149054 263640 150484
rect 263600 149048 263652 149054
rect 263600 148990 263652 148996
rect 262864 148844 262916 148850
rect 262864 148786 262916 148792
rect 262588 147756 262640 147762
rect 262588 147698 262640 147704
rect 260932 3596 260984 3602
rect 260932 3538 260984 3544
rect 262876 3534 262904 148786
rect 263508 148776 263560 148782
rect 263508 148718 263560 148724
rect 263520 3534 263548 148718
rect 264256 148306 264284 150484
rect 264624 150470 264914 150498
rect 264244 148300 264296 148306
rect 264244 148242 264296 148248
rect 264624 148170 264652 150470
rect 264888 148912 264940 148918
rect 264888 148854 264940 148860
rect 264612 148164 264664 148170
rect 264612 148106 264664 148112
rect 264900 3534 264928 148854
rect 265636 148374 265664 150484
rect 265624 148368 265676 148374
rect 265624 148310 265676 148316
rect 266280 147830 266308 150484
rect 267016 148238 267044 150484
rect 267108 150470 267674 150498
rect 267004 148232 267056 148238
rect 267004 148174 267056 148180
rect 266268 147824 266320 147830
rect 266268 147766 266320 147772
rect 267108 146282 267136 150470
rect 268396 148442 268424 150484
rect 268672 150470 269054 150498
rect 268384 148436 268436 148442
rect 268384 148378 268436 148384
rect 267188 148368 267240 148374
rect 267188 148310 267240 148316
rect 266464 146254 267136 146282
rect 266464 3670 266492 146254
rect 267200 142154 267228 148310
rect 267648 148232 267700 148238
rect 267648 148174 267700 148180
rect 267016 142126 267228 142154
rect 266452 3664 266504 3670
rect 266452 3606 266504 3612
rect 267016 3534 267044 142126
rect 260748 3528 260800 3534
rect 260748 3470 260800 3476
rect 261760 3528 261812 3534
rect 261760 3470 261812 3476
rect 262864 3528 262916 3534
rect 262864 3470 262916 3476
rect 262956 3528 263008 3534
rect 262956 3470 263008 3476
rect 263508 3528 263560 3534
rect 263508 3470 263560 3476
rect 264152 3528 264204 3534
rect 264152 3470 264204 3476
rect 264888 3528 264940 3534
rect 264888 3470 264940 3476
rect 265348 3528 265400 3534
rect 265348 3470 265400 3476
rect 267004 3528 267056 3534
rect 267004 3470 267056 3476
rect 261772 480 261800 3470
rect 262968 480 262996 3470
rect 264164 480 264192 3470
rect 265360 480 265388 3470
rect 267660 3194 267688 148174
rect 268672 148034 268700 150470
rect 268936 148436 268988 148442
rect 268936 148378 268988 148384
rect 268660 148028 268712 148034
rect 268660 147970 268712 147976
rect 268948 3602 268976 148378
rect 269028 148300 269080 148306
rect 269028 148242 269080 148248
rect 267740 3596 267792 3602
rect 267740 3538 267792 3544
rect 268936 3596 268988 3602
rect 268936 3538 268988 3544
rect 266544 3188 266596 3194
rect 266544 3130 266596 3136
rect 267648 3188 267700 3194
rect 267648 3130 267700 3136
rect 266556 480 266584 3130
rect 267752 480 267780 3538
rect 269040 3482 269068 148242
rect 269776 148102 269804 150484
rect 269868 150470 270434 150498
rect 269764 148096 269816 148102
rect 269764 148038 269816 148044
rect 269868 142154 269896 150470
rect 270408 149048 270460 149054
rect 270408 148990 270460 148996
rect 269224 142126 269896 142154
rect 269224 3738 269252 142126
rect 269212 3732 269264 3738
rect 269212 3674 269264 3680
rect 268856 3454 269068 3482
rect 268856 480 268884 3454
rect 270052 598 270264 626
rect 270052 480 270080 598
rect 270236 490 270264 598
rect 270420 490 270448 148990
rect 271156 148578 271184 150484
rect 271432 150470 271814 150498
rect 271144 148572 271196 148578
rect 271144 148514 271196 148520
rect 271432 147966 271460 150470
rect 271788 148572 271840 148578
rect 271788 148514 271840 148520
rect 271420 147960 271472 147966
rect 271420 147902 271472 147908
rect 271800 3330 271828 148514
rect 272536 148510 272564 150484
rect 272524 148504 272576 148510
rect 272524 148446 272576 148452
rect 273180 147898 273208 150484
rect 273824 148714 273852 150484
rect 274560 148986 274588 150484
rect 274548 148980 274600 148986
rect 274548 148922 274600 148928
rect 273812 148708 273864 148714
rect 273812 148650 273864 148656
rect 274548 148708 274600 148714
rect 274548 148650 274600 148656
rect 273904 148504 273956 148510
rect 273904 148446 273956 148452
rect 273168 147892 273220 147898
rect 273168 147834 273220 147840
rect 273628 3528 273680 3534
rect 273628 3470 273680 3476
rect 272432 3460 272484 3466
rect 272432 3402 272484 3408
rect 271236 3324 271288 3330
rect 271236 3266 271288 3272
rect 271788 3324 271840 3330
rect 271788 3266 271840 3272
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270236 462 270448 490
rect 271248 480 271276 3266
rect 272444 480 272472 3402
rect 273640 480 273668 3470
rect 273916 3466 273944 148446
rect 274560 3534 274588 148650
rect 275204 148646 275232 150484
rect 275940 148850 275968 150484
rect 275928 148844 275980 148850
rect 275928 148786 275980 148792
rect 276584 148782 276612 150484
rect 276952 150470 277334 150498
rect 276952 148918 276980 150470
rect 276940 148912 276992 148918
rect 276940 148854 276992 148860
rect 277216 148912 277268 148918
rect 277216 148854 277268 148860
rect 276572 148776 276624 148782
rect 276572 148718 276624 148724
rect 276664 148776 276716 148782
rect 276664 148718 276716 148724
rect 275192 148640 275244 148646
rect 275192 148582 275244 148588
rect 276020 3596 276072 3602
rect 276020 3538 276072 3544
rect 274548 3528 274600 3534
rect 274548 3470 274600 3476
rect 273904 3460 273956 3466
rect 273904 3402 273956 3408
rect 274824 3052 274876 3058
rect 274824 2994 274876 3000
rect 274836 480 274864 2994
rect 276032 480 276060 3538
rect 276676 3058 276704 148718
rect 277228 3602 277256 148854
rect 277308 148640 277360 148646
rect 277308 148582 277360 148588
rect 277216 3596 277268 3602
rect 277216 3538 277268 3544
rect 277320 3482 277348 148582
rect 277964 148374 277992 150484
rect 277952 148368 278004 148374
rect 277952 148310 278004 148316
rect 278700 148238 278728 150484
rect 279344 148442 279372 150484
rect 279332 148436 279384 148442
rect 279332 148378 279384 148384
rect 280080 148306 280108 150484
rect 280724 149054 280752 150484
rect 280712 149048 280764 149054
rect 280712 148990 280764 148996
rect 281368 148578 281396 150484
rect 281356 148572 281408 148578
rect 281356 148514 281408 148520
rect 282104 148510 282132 150484
rect 282748 148714 282776 150484
rect 283484 148782 283512 150484
rect 284128 148918 284156 150484
rect 284116 148912 284168 148918
rect 284116 148854 284168 148860
rect 283472 148776 283524 148782
rect 283472 148718 283524 148724
rect 282736 148708 282788 148714
rect 282736 148650 282788 148656
rect 284864 148646 284892 150484
rect 284852 148640 284904 148646
rect 284852 148582 284904 148588
rect 282092 148504 282144 148510
rect 282092 148446 282144 148452
rect 280068 148300 280120 148306
rect 280068 148242 280120 148248
rect 278688 148232 278740 148238
rect 278688 148174 278740 148180
rect 285508 148034 285536 150484
rect 278688 148028 278740 148034
rect 278688 147970 278740 147976
rect 285496 148028 285548 148034
rect 285496 147970 285548 147976
rect 277136 3454 277348 3482
rect 276664 3052 276716 3058
rect 276664 2994 276716 3000
rect 277136 480 277164 3454
rect 278332 598 278544 626
rect 278332 480 278360 598
rect 278516 490 278544 598
rect 278700 490 278728 147970
rect 286244 147966 286272 150484
rect 280804 147960 280856 147966
rect 280804 147902 280856 147908
rect 286232 147960 286284 147966
rect 286232 147902 286284 147908
rect 280712 3528 280764 3534
rect 280712 3470 280764 3476
rect 279516 3460 279568 3466
rect 279516 3402 279568 3408
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 278516 462 278728 490
rect 279528 480 279556 3402
rect 280724 480 280752 3470
rect 280816 3466 280844 147902
rect 286888 147898 286916 150484
rect 286968 148436 287020 148442
rect 286968 148378 287020 148384
rect 281448 147892 281500 147898
rect 281448 147834 281500 147840
rect 286876 147892 286928 147898
rect 286876 147834 286928 147840
rect 281460 3534 281488 147834
rect 282828 147824 282880 147830
rect 282828 147766 282880 147772
rect 281448 3528 281500 3534
rect 281448 3470 281500 3476
rect 280804 3460 280856 3466
rect 280804 3402 280856 3408
rect 282840 3058 282868 147766
rect 285496 147756 285548 147762
rect 285496 147698 285548 147704
rect 285508 6914 285536 147698
rect 285588 147688 285640 147694
rect 285588 147630 285640 147636
rect 285416 6886 285536 6914
rect 283104 3800 283156 3806
rect 283104 3742 283156 3748
rect 281908 3052 281960 3058
rect 281908 2994 281960 3000
rect 282828 3052 282880 3058
rect 282828 2994 282880 3000
rect 281920 480 281948 2994
rect 283116 480 283144 3742
rect 284300 3528 284352 3534
rect 284300 3470 284352 3476
rect 284312 480 284340 3470
rect 285416 480 285444 6886
rect 285600 3534 285628 147630
rect 285588 3528 285640 3534
rect 285588 3470 285640 3476
rect 286612 598 286824 626
rect 286612 480 286640 598
rect 286796 490 286824 598
rect 286980 490 287008 148378
rect 287624 147830 287652 150484
rect 287900 150470 288282 150498
rect 287612 147824 287664 147830
rect 287612 147766 287664 147772
rect 287900 142154 287928 150470
rect 288348 147756 288400 147762
rect 288348 147698 288400 147704
rect 287164 142126 287928 142154
rect 287164 3806 287192 142126
rect 287152 3800 287204 3806
rect 287152 3742 287204 3748
rect 288360 3534 288388 147698
rect 289004 147694 289032 150484
rect 289648 147830 289676 150484
rect 290292 148442 290320 150484
rect 290280 148436 290332 148442
rect 290280 148378 290332 148384
rect 289636 147824 289688 147830
rect 289636 147766 289688 147772
rect 291028 147762 291056 150484
rect 291016 147756 291068 147762
rect 291016 147698 291068 147704
rect 291672 147694 291700 150484
rect 291764 150470 292422 150498
rect 292592 150470 293066 150498
rect 293236 150470 293802 150498
rect 293972 150470 294446 150498
rect 294616 150470 295182 150498
rect 295444 150470 295826 150498
rect 296562 150470 296668 150498
rect 288992 147688 289044 147694
rect 288992 147630 289044 147636
rect 289728 147688 289780 147694
rect 289728 147630 289780 147636
rect 291660 147688 291712 147694
rect 291660 147630 291712 147636
rect 289740 3534 289768 147630
rect 291764 142154 291792 150470
rect 292592 147778 292620 150470
rect 291304 142126 291792 142154
rect 292500 147750 292620 147778
rect 291304 3534 291332 142126
rect 292500 3534 292528 147750
rect 293236 142154 293264 150470
rect 292776 142126 293264 142154
rect 292776 6914 292804 142126
rect 292592 6886 292804 6914
rect 287796 3528 287848 3534
rect 287796 3470 287848 3476
rect 288348 3528 288400 3534
rect 288348 3470 288400 3476
rect 288992 3528 289044 3534
rect 288992 3470 289044 3476
rect 289728 3528 289780 3534
rect 289728 3470 289780 3476
rect 290188 3528 290240 3534
rect 290188 3470 290240 3476
rect 291292 3528 291344 3534
rect 291292 3470 291344 3476
rect 291384 3528 291436 3534
rect 291384 3470 291436 3476
rect 292488 3528 292540 3534
rect 292488 3470 292540 3476
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 286796 462 287008 490
rect 287808 480 287836 3470
rect 289004 480 289032 3470
rect 290200 480 290228 3470
rect 291396 480 291424 3470
rect 292592 480 292620 6886
rect 293972 2802 294000 150470
rect 294616 142154 294644 150470
rect 294064 142126 294644 142154
rect 294064 3534 294092 142126
rect 295444 3534 295472 150470
rect 296640 4146 296668 150470
rect 297192 147694 297220 150484
rect 297836 147762 297864 150484
rect 297824 147756 297876 147762
rect 297824 147698 297876 147704
rect 298572 147694 298600 150484
rect 299230 150470 299428 150498
rect 298744 147756 298796 147762
rect 298744 147698 298796 147704
rect 297180 147688 297232 147694
rect 297180 147630 297232 147636
rect 298284 147688 298336 147694
rect 298284 147630 298336 147636
rect 298560 147688 298612 147694
rect 298560 147630 298612 147636
rect 298296 16574 298324 147630
rect 298296 16546 298508 16574
rect 296628 4140 296680 4146
rect 296628 4082 296680 4088
rect 297272 4140 297324 4146
rect 297272 4082 297324 4088
rect 294052 3528 294104 3534
rect 294052 3470 294104 3476
rect 294880 3528 294932 3534
rect 294880 3470 294932 3476
rect 295432 3528 295484 3534
rect 295432 3470 295484 3476
rect 296076 3528 296128 3534
rect 296076 3470 296128 3476
rect 293696 2774 294000 2802
rect 293696 480 293724 2774
rect 294892 480 294920 3470
rect 296088 480 296116 3470
rect 297284 480 297312 4082
rect 298480 480 298508 16546
rect 298756 3534 298784 147698
rect 298744 3528 298796 3534
rect 298744 3470 298796 3476
rect 299400 3126 299428 150470
rect 299952 147694 299980 150484
rect 300610 150470 300808 150498
rect 299664 147688 299716 147694
rect 299664 147630 299716 147636
rect 299940 147688 299992 147694
rect 299940 147630 299992 147636
rect 299676 16574 299704 147630
rect 299676 16546 300716 16574
rect 299664 3528 299716 3534
rect 299664 3470 299716 3476
rect 299388 3120 299440 3126
rect 299388 3062 299440 3068
rect 299676 480 299704 3470
rect 300688 3210 300716 16546
rect 300780 3330 300808 150470
rect 301332 147762 301360 150484
rect 301976 147830 302004 150484
rect 301964 147824 302016 147830
rect 301964 147766 302016 147772
rect 301320 147756 301372 147762
rect 301320 147698 301372 147704
rect 302712 147694 302740 150484
rect 303370 150470 303568 150498
rect 304106 150470 304580 150498
rect 304750 150470 304948 150498
rect 302424 147688 302476 147694
rect 302424 147630 302476 147636
rect 302700 147688 302752 147694
rect 302700 147630 302752 147636
rect 303436 147688 303488 147694
rect 303436 147630 303488 147636
rect 302436 16574 302464 147630
rect 302436 16546 303200 16574
rect 300768 3324 300820 3330
rect 300768 3266 300820 3272
rect 300688 3182 300808 3210
rect 300780 480 300808 3182
rect 301964 3120 302016 3126
rect 301964 3062 302016 3068
rect 301976 480 302004 3062
rect 303172 480 303200 16546
rect 303448 2990 303476 147630
rect 303540 4146 303568 150470
rect 304552 142154 304580 150470
rect 304552 142126 304856 142154
rect 303528 4140 303580 4146
rect 303528 4082 303580 4088
rect 304828 3806 304856 142126
rect 304816 3800 304868 3806
rect 304816 3742 304868 3748
rect 304920 3670 304948 150470
rect 305184 147756 305236 147762
rect 305184 147698 305236 147704
rect 305196 16574 305224 147698
rect 305472 147694 305500 150484
rect 306130 150470 306328 150498
rect 305460 147688 305512 147694
rect 305460 147630 305512 147636
rect 306196 147688 306248 147694
rect 306196 147630 306248 147636
rect 305196 16546 305592 16574
rect 304908 3664 304960 3670
rect 304908 3606 304960 3612
rect 304356 3324 304408 3330
rect 304356 3266 304408 3272
rect 303436 2984 303488 2990
rect 303436 2926 303488 2932
rect 304368 480 304396 3266
rect 305564 480 305592 16546
rect 306208 3602 306236 147630
rect 306196 3596 306248 3602
rect 306196 3538 306248 3544
rect 306300 3466 306328 150470
rect 306564 147824 306616 147830
rect 306564 147766 306616 147772
rect 306576 16574 306604 147766
rect 306760 147694 306788 150484
rect 307510 150470 307616 150498
rect 306748 147688 306800 147694
rect 306748 147630 306800 147636
rect 306576 16546 306788 16574
rect 306288 3460 306340 3466
rect 306288 3402 306340 3408
rect 306760 480 306788 16546
rect 307588 4010 307616 150470
rect 308140 147694 308168 150484
rect 308876 147830 308904 150484
rect 308864 147824 308916 147830
rect 308864 147766 308916 147772
rect 309520 147762 309548 150484
rect 310270 150470 310376 150498
rect 309508 147756 309560 147762
rect 309508 147698 309560 147704
rect 307668 147688 307720 147694
rect 307668 147630 307720 147636
rect 308128 147688 308180 147694
rect 308128 147630 308180 147636
rect 309784 147688 309836 147694
rect 309784 147630 309836 147636
rect 307576 4004 307628 4010
rect 307576 3946 307628 3952
rect 307680 3534 307708 147630
rect 309048 4140 309100 4146
rect 309048 4082 309100 4088
rect 307668 3528 307720 3534
rect 307668 3470 307720 3476
rect 307944 2984 307996 2990
rect 307944 2926 307996 2932
rect 307956 480 307984 2926
rect 309060 480 309088 4082
rect 309796 3874 309824 147630
rect 309784 3868 309836 3874
rect 309784 3810 309836 3816
rect 310244 3800 310296 3806
rect 310244 3742 310296 3748
rect 310256 480 310284 3742
rect 310348 3738 310376 150470
rect 310428 147756 310480 147762
rect 310428 147698 310480 147704
rect 310440 3942 310468 147698
rect 310900 147694 310928 150484
rect 311636 148374 311664 150484
rect 311624 148368 311676 148374
rect 311624 148310 311676 148316
rect 311164 147824 311216 147830
rect 311164 147766 311216 147772
rect 310888 147688 310940 147694
rect 310888 147630 310940 147636
rect 310428 3936 310480 3942
rect 310428 3878 310480 3884
rect 310336 3732 310388 3738
rect 310336 3674 310388 3680
rect 311176 3262 311204 147766
rect 312280 147694 312308 150484
rect 313016 147762 313044 150484
rect 313004 147756 313056 147762
rect 313004 147698 313056 147704
rect 313660 147694 313688 150484
rect 314318 150470 314608 150498
rect 313924 147756 313976 147762
rect 313924 147698 313976 147704
rect 311808 147688 311860 147694
rect 311808 147630 311860 147636
rect 312268 147688 312320 147694
rect 312268 147630 312320 147636
rect 313188 147688 313240 147694
rect 313188 147630 313240 147636
rect 313648 147688 313700 147694
rect 313648 147630 313700 147636
rect 311820 3806 311848 147630
rect 311808 3800 311860 3806
rect 311808 3742 311860 3748
rect 313200 3670 313228 147630
rect 311440 3664 311492 3670
rect 311440 3606 311492 3612
rect 313188 3664 313240 3670
rect 313188 3606 313240 3612
rect 311164 3256 311216 3262
rect 311164 3198 311216 3204
rect 311452 480 311480 3606
rect 312636 3596 312688 3602
rect 312636 3538 312688 3544
rect 312648 480 312676 3538
rect 313832 3460 313884 3466
rect 313832 3402 313884 3408
rect 313844 480 313872 3402
rect 313936 3398 313964 147698
rect 314476 147688 314528 147694
rect 314476 147630 314528 147636
rect 314488 3466 314516 147630
rect 314580 3602 314608 150470
rect 315040 147762 315068 150484
rect 315698 150470 315988 150498
rect 315028 147756 315080 147762
rect 315028 147698 315080 147704
rect 315960 4146 315988 150470
rect 316420 147694 316448 150484
rect 317078 150470 317368 150498
rect 316408 147688 316460 147694
rect 316408 147630 316460 147636
rect 317236 147688 317288 147694
rect 317236 147630 317288 147636
rect 315948 4140 316000 4146
rect 315948 4082 316000 4088
rect 317248 4078 317276 147630
rect 317236 4072 317288 4078
rect 317236 4014 317288 4020
rect 317340 4026 317368 150470
rect 317800 147694 317828 150484
rect 318458 150470 318748 150498
rect 318064 147756 318116 147762
rect 318064 147698 318116 147704
rect 317788 147688 317840 147694
rect 317788 147630 317840 147636
rect 317340 3998 317460 4026
rect 317432 3874 317460 3998
rect 317328 3868 317380 3874
rect 317328 3810 317380 3816
rect 317420 3868 317472 3874
rect 317420 3810 317472 3816
rect 316224 3732 316276 3738
rect 316224 3674 316276 3680
rect 314568 3596 314620 3602
rect 314568 3538 314620 3544
rect 315028 3528 315080 3534
rect 315028 3470 315080 3476
rect 314476 3460 314528 3466
rect 314476 3402 314528 3408
rect 313924 3392 313976 3398
rect 313924 3334 313976 3340
rect 315040 480 315068 3470
rect 316236 480 316264 3674
rect 317340 480 317368 3810
rect 318076 3330 318104 147698
rect 318616 147688 318668 147694
rect 318616 147630 318668 147636
rect 318064 3324 318116 3330
rect 318064 3266 318116 3272
rect 318524 3256 318576 3262
rect 318524 3198 318576 3204
rect 318536 480 318564 3198
rect 318628 2990 318656 147630
rect 318720 4010 318748 150470
rect 319180 147694 319208 150484
rect 319838 150470 320036 150498
rect 319168 147688 319220 147694
rect 319168 147630 319220 147636
rect 318708 4004 318760 4010
rect 318708 3946 318760 3952
rect 319720 3936 319772 3942
rect 319720 3878 319772 3884
rect 318616 2984 318668 2990
rect 318616 2926 318668 2932
rect 319732 480 319760 3878
rect 320008 3874 320036 150470
rect 320560 147694 320588 150484
rect 321218 150470 321508 150498
rect 320088 147688 320140 147694
rect 320088 147630 320140 147636
rect 320548 147688 320600 147694
rect 320548 147630 320600 147636
rect 321376 147688 321428 147694
rect 321376 147630 321428 147636
rect 319996 3868 320048 3874
rect 319996 3810 320048 3816
rect 320100 3058 320128 147630
rect 321388 4826 321416 147630
rect 321376 4820 321428 4826
rect 321376 4762 321428 4768
rect 321480 3738 321508 150470
rect 321940 147694 321968 150484
rect 322584 148510 322612 150484
rect 322572 148504 322624 148510
rect 322572 148446 322624 148452
rect 322204 148368 322256 148374
rect 322204 148310 322256 148316
rect 321928 147688 321980 147694
rect 321928 147630 321980 147636
rect 322112 3800 322164 3806
rect 322112 3742 322164 3748
rect 321468 3732 321520 3738
rect 321468 3674 321520 3680
rect 320916 3528 320968 3534
rect 320916 3470 320968 3476
rect 320088 3052 320140 3058
rect 320088 2994 320140 3000
rect 320928 480 320956 3470
rect 322124 480 322152 3742
rect 322216 3534 322244 148310
rect 323228 147694 323256 150484
rect 323978 150470 324176 150498
rect 322848 147688 322900 147694
rect 322848 147630 322900 147636
rect 323216 147688 323268 147694
rect 323216 147630 323268 147636
rect 322860 3806 322888 147630
rect 322848 3800 322900 3806
rect 322848 3742 322900 3748
rect 324148 3534 324176 150470
rect 324608 147694 324636 150484
rect 325358 150470 325648 150498
rect 324228 147688 324280 147694
rect 324228 147630 324280 147636
rect 324596 147688 324648 147694
rect 324596 147630 324648 147636
rect 325516 147688 325568 147694
rect 325516 147630 325568 147636
rect 322204 3528 322256 3534
rect 322204 3470 322256 3476
rect 323308 3528 323360 3534
rect 323308 3470 323360 3476
rect 324136 3528 324188 3534
rect 324136 3470 324188 3476
rect 323320 480 323348 3470
rect 324240 3126 324268 147630
rect 325528 5166 325556 147630
rect 325516 5160 325568 5166
rect 325516 5102 325568 5108
rect 325620 3670 325648 150470
rect 325988 147694 326016 150484
rect 326724 148442 326752 150484
rect 326712 148436 326764 148442
rect 326712 148378 326764 148384
rect 327368 147694 327396 150484
rect 328118 150470 328408 150498
rect 325976 147688 326028 147694
rect 325976 147630 326028 147636
rect 326988 147688 327040 147694
rect 326988 147630 327040 147636
rect 327356 147688 327408 147694
rect 327356 147630 327408 147636
rect 328276 147688 328328 147694
rect 328276 147630 328328 147636
rect 324412 3664 324464 3670
rect 324412 3606 324464 3612
rect 325608 3664 325660 3670
rect 325608 3606 325660 3612
rect 324228 3120 324280 3126
rect 324228 3062 324280 3068
rect 324424 480 324452 3606
rect 327000 3466 327028 147630
rect 328000 3596 328052 3602
rect 328000 3538 328052 3544
rect 326804 3460 326856 3466
rect 326804 3402 326856 3408
rect 326988 3460 327040 3466
rect 326988 3402 327040 3408
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 325620 480 325648 3334
rect 326816 480 326844 3402
rect 328012 480 328040 3538
rect 328288 3194 328316 147630
rect 328380 3602 328408 150470
rect 328748 148578 328776 150484
rect 329498 150470 329788 150498
rect 328736 148572 328788 148578
rect 328736 148514 328788 148520
rect 328368 3596 328420 3602
rect 328368 3538 328420 3544
rect 329760 3330 329788 150470
rect 330128 147694 330156 150484
rect 330772 148374 330800 150484
rect 330760 148368 330812 148374
rect 330760 148310 330812 148316
rect 331508 147694 331536 150484
rect 332166 150470 332548 150498
rect 330116 147688 330168 147694
rect 330116 147630 330168 147636
rect 331128 147688 331180 147694
rect 331128 147630 331180 147636
rect 331496 147688 331548 147694
rect 331496 147630 331548 147636
rect 332416 147688 332468 147694
rect 332416 147630 332468 147636
rect 330392 4140 330444 4146
rect 330392 4082 330444 4088
rect 329196 3324 329248 3330
rect 329196 3266 329248 3272
rect 329748 3324 329800 3330
rect 329748 3266 329800 3272
rect 328276 3188 328328 3194
rect 328276 3130 328328 3136
rect 329208 480 329236 3266
rect 330404 480 330432 4082
rect 331140 3262 331168 147630
rect 332428 4146 332456 147630
rect 332416 4140 332468 4146
rect 332416 4082 332468 4088
rect 331588 4072 331640 4078
rect 331588 4014 331640 4020
rect 331128 3256 331180 3262
rect 331128 3198 331180 3204
rect 331600 480 331628 4014
rect 332520 3398 332548 150470
rect 332888 147762 332916 150484
rect 333546 150470 333928 150498
rect 332876 147756 332928 147762
rect 332876 147698 332928 147704
rect 333900 4078 333928 150470
rect 334268 147694 334296 150484
rect 334926 150470 335216 150498
rect 334624 147756 334676 147762
rect 334624 147698 334676 147704
rect 334256 147688 334308 147694
rect 334256 147630 334308 147636
rect 334636 7682 334664 147698
rect 334624 7676 334676 7682
rect 334624 7618 334676 7624
rect 335188 4894 335216 150470
rect 335648 147694 335676 150484
rect 336306 150470 336688 150498
rect 335268 147688 335320 147694
rect 335268 147630 335320 147636
rect 335636 147688 335688 147694
rect 335636 147630 335688 147636
rect 336556 147688 336608 147694
rect 336556 147630 336608 147636
rect 335176 4888 335228 4894
rect 335176 4830 335228 4836
rect 333888 4072 333940 4078
rect 333888 4014 333940 4020
rect 335280 4010 335308 147630
rect 336568 4962 336596 147630
rect 336556 4956 336608 4962
rect 336556 4898 336608 4904
rect 332692 4004 332744 4010
rect 332692 3946 332744 3952
rect 335268 4004 335320 4010
rect 335268 3946 335320 3952
rect 332508 3392 332560 3398
rect 332508 3334 332560 3340
rect 332704 480 332732 3946
rect 336660 3942 336688 150470
rect 337028 147762 337056 150484
rect 337672 147830 337700 150484
rect 337660 147824 337712 147830
rect 337660 147766 337712 147772
rect 337016 147756 337068 147762
rect 337016 147698 337068 147704
rect 338408 147694 338436 150484
rect 339066 150470 339356 150498
rect 338764 148504 338816 148510
rect 338764 148446 338816 148452
rect 338396 147688 338448 147694
rect 338396 147630 338448 147636
rect 338672 4820 338724 4826
rect 338672 4762 338724 4768
rect 335084 3936 335136 3942
rect 335084 3878 335136 3884
rect 336648 3936 336700 3942
rect 336648 3878 336700 3884
rect 333888 2984 333940 2990
rect 333888 2926 333940 2932
rect 333900 480 333928 2926
rect 335096 480 335124 3878
rect 337476 3868 337528 3874
rect 337476 3810 337528 3816
rect 336280 3052 336332 3058
rect 336280 2994 336332 3000
rect 336292 480 336320 2994
rect 337488 480 337516 3810
rect 338684 480 338712 4762
rect 338776 4214 338804 148446
rect 339328 15910 339356 150470
rect 339696 147694 339724 150484
rect 340446 150470 340828 150498
rect 340144 147756 340196 147762
rect 340144 147698 340196 147704
rect 339408 147688 339460 147694
rect 339408 147630 339460 147636
rect 339684 147688 339736 147694
rect 339684 147630 339736 147636
rect 339316 15904 339368 15910
rect 339316 15846 339368 15852
rect 338764 4208 338816 4214
rect 338764 4150 338816 4156
rect 339420 3874 339448 147630
rect 340156 5030 340184 147698
rect 340696 147688 340748 147694
rect 340696 147630 340748 147636
rect 340708 18630 340736 147630
rect 340696 18624 340748 18630
rect 340696 18566 340748 18572
rect 340144 5024 340196 5030
rect 340144 4966 340196 4972
rect 339408 3868 339460 3874
rect 339408 3810 339460 3816
rect 340800 3738 340828 150470
rect 341076 147694 341104 150484
rect 341826 150470 342116 150498
rect 341064 147688 341116 147694
rect 341064 147630 341116 147636
rect 342088 6594 342116 150470
rect 342456 147694 342484 150484
rect 343206 150470 343496 150498
rect 342904 147824 342956 147830
rect 342904 147766 342956 147772
rect 342168 147688 342220 147694
rect 342168 147630 342220 147636
rect 342444 147688 342496 147694
rect 342444 147630 342496 147636
rect 342076 6588 342128 6594
rect 342076 6530 342128 6536
rect 342180 4826 342208 147630
rect 342916 5098 342944 147766
rect 343468 8974 343496 150470
rect 343836 147762 343864 150484
rect 344586 150470 344968 150498
rect 343824 147756 343876 147762
rect 343824 147698 343876 147704
rect 343548 147688 343600 147694
rect 343548 147630 343600 147636
rect 343456 8968 343508 8974
rect 343456 8910 343508 8916
rect 342904 5092 342956 5098
rect 342904 5034 342956 5040
rect 342168 4820 342220 4826
rect 342168 4762 342220 4768
rect 342168 4208 342220 4214
rect 342168 4150 342220 4156
rect 340972 3800 341024 3806
rect 340972 3742 341024 3748
rect 339868 3732 339920 3738
rect 339868 3674 339920 3680
rect 340788 3732 340840 3738
rect 340788 3674 340840 3680
rect 339880 480 339908 3674
rect 340984 480 341012 3742
rect 342180 480 342208 4150
rect 343560 3806 343588 147630
rect 343548 3800 343600 3806
rect 343548 3742 343600 3748
rect 344940 3534 344968 150470
rect 345216 147694 345244 150484
rect 345966 150470 346348 150498
rect 345664 147756 345716 147762
rect 345664 147698 345716 147704
rect 345204 147688 345256 147694
rect 345204 147630 345256 147636
rect 345676 25566 345704 147698
rect 346216 147688 346268 147694
rect 346216 147630 346268 147636
rect 345664 25560 345716 25566
rect 345664 25502 345716 25508
rect 346228 6526 346256 147630
rect 346216 6520 346268 6526
rect 346216 6462 346268 6468
rect 346320 6458 346348 150470
rect 346596 147694 346624 150484
rect 347240 148510 347268 150484
rect 347976 148986 348004 150484
rect 348634 150470 349108 150498
rect 347964 148980 348016 148986
rect 347964 148922 348016 148928
rect 347228 148504 347280 148510
rect 347228 148446 347280 148452
rect 346584 147688 346636 147694
rect 346584 147630 346636 147636
rect 347688 147688 347740 147694
rect 347688 147630 347740 147636
rect 346308 6452 346360 6458
rect 346308 6394 346360 6400
rect 345756 5160 345808 5166
rect 345756 5102 345808 5108
rect 344560 3528 344612 3534
rect 344560 3470 344612 3476
rect 344928 3528 344980 3534
rect 344928 3470 344980 3476
rect 343364 3120 343416 3126
rect 343364 3062 343416 3068
rect 343376 480 343404 3062
rect 344572 480 344600 3470
rect 345768 480 345796 5102
rect 347700 3670 347728 147630
rect 346952 3664 347004 3670
rect 346952 3606 347004 3612
rect 347688 3664 347740 3670
rect 347688 3606 347740 3612
rect 346964 480 346992 3606
rect 349080 3466 349108 150470
rect 349356 148918 349384 150484
rect 350014 150470 350488 150498
rect 349344 148912 349396 148918
rect 349344 148854 349396 148860
rect 349252 148436 349304 148442
rect 349252 148378 349304 148384
rect 348056 3460 348108 3466
rect 348056 3402 348108 3408
rect 349068 3460 349120 3466
rect 349068 3402 349120 3408
rect 348068 480 348096 3402
rect 349264 480 349292 148378
rect 350460 6390 350488 150470
rect 350736 147694 350764 150484
rect 351380 148850 351408 150484
rect 351368 148844 351420 148850
rect 351368 148786 351420 148792
rect 352012 148572 352064 148578
rect 352012 148514 352064 148520
rect 350724 147688 350776 147694
rect 350724 147630 350776 147636
rect 351828 147688 351880 147694
rect 351828 147630 351880 147636
rect 350448 6384 350500 6390
rect 350448 6326 350500 6332
rect 351840 3602 351868 147630
rect 352024 16574 352052 148514
rect 352116 147694 352144 150484
rect 352760 148782 352788 150484
rect 352748 148776 352800 148782
rect 352748 148718 352800 148724
rect 353496 147694 353524 150484
rect 354154 150470 354536 150498
rect 352104 147688 352156 147694
rect 352104 147630 352156 147636
rect 353208 147688 353260 147694
rect 353208 147630 353260 147636
rect 353484 147688 353536 147694
rect 353484 147630 353536 147636
rect 352024 16546 352880 16574
rect 351644 3596 351696 3602
rect 351644 3538 351696 3544
rect 351828 3596 351880 3602
rect 351828 3538 351880 3544
rect 350448 3188 350500 3194
rect 350448 3130 350500 3136
rect 350460 480 350488 3130
rect 351656 480 351684 3538
rect 352852 480 352880 16546
rect 353220 6322 353248 147630
rect 353208 6316 353260 6322
rect 353208 6258 353260 6264
rect 354508 6186 354536 150470
rect 354876 147694 354904 150484
rect 355534 150470 355916 150498
rect 354588 147688 354640 147694
rect 354588 147630 354640 147636
rect 354864 147688 354916 147694
rect 354864 147630 354916 147636
rect 354496 6180 354548 6186
rect 354496 6122 354548 6128
rect 354600 4282 354628 147630
rect 355888 4418 355916 150470
rect 356164 148578 356192 150484
rect 356900 148714 356928 150484
rect 356888 148708 356940 148714
rect 356888 148650 356940 148656
rect 356152 148572 356204 148578
rect 356152 148514 356204 148520
rect 357348 148572 357400 148578
rect 357348 148514 357400 148520
rect 356152 148368 356204 148374
rect 356152 148310 356204 148316
rect 355968 147688 356020 147694
rect 355968 147630 356020 147636
rect 355876 4412 355928 4418
rect 355876 4354 355928 4360
rect 354588 4276 354640 4282
rect 354588 4218 354640 4224
rect 354036 3324 354088 3330
rect 354036 3266 354088 3272
rect 354048 480 354076 3266
rect 355232 3256 355284 3262
rect 355232 3198 355284 3204
rect 355244 480 355272 3198
rect 355980 3126 356008 147630
rect 356164 16574 356192 148310
rect 356164 16546 356376 16574
rect 355968 3120 356020 3126
rect 355968 3062 356020 3068
rect 356348 480 356376 16546
rect 357360 6254 357388 148514
rect 357544 147694 357572 150484
rect 358294 150470 358676 150498
rect 357532 147688 357584 147694
rect 357532 147630 357584 147636
rect 358648 7614 358676 150470
rect 358924 147694 358952 150484
rect 359674 150470 360056 150498
rect 358728 147688 358780 147694
rect 358728 147630 358780 147636
rect 358912 147688 358964 147694
rect 358912 147630 358964 147636
rect 358636 7608 358688 7614
rect 358636 7550 358688 7556
rect 357348 6248 357400 6254
rect 357348 6190 357400 6196
rect 358740 4350 358768 147630
rect 359924 7676 359976 7682
rect 359924 7618 359976 7624
rect 358728 4344 358780 4350
rect 358728 4286 358780 4292
rect 357532 4140 357584 4146
rect 357532 4082 357584 4088
rect 357544 480 357572 4082
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 359936 480 359964 7618
rect 360028 4554 360056 150470
rect 360304 148578 360332 150484
rect 361054 150470 361528 150498
rect 360292 148572 360344 148578
rect 360292 148514 360344 148520
rect 360108 147688 360160 147694
rect 360108 147630 360160 147636
rect 360016 4548 360068 4554
rect 360016 4490 360068 4496
rect 360120 3194 360148 147630
rect 361120 4072 361172 4078
rect 361120 4014 361172 4020
rect 360108 3188 360160 3194
rect 360108 3130 360160 3136
rect 361132 480 361160 4014
rect 361500 3262 361528 150470
rect 361684 147694 361712 150484
rect 362434 150470 362908 150498
rect 362880 147778 362908 150470
rect 362880 147750 363000 147778
rect 361672 147688 361724 147694
rect 361672 147630 361724 147636
rect 362868 147688 362920 147694
rect 362868 147630 362920 147636
rect 362880 4486 362908 147630
rect 362972 147082 363000 147750
rect 363064 147694 363092 150484
rect 363722 150470 364196 150498
rect 363052 147688 363104 147694
rect 363052 147630 363104 147636
rect 362960 147076 363012 147082
rect 362960 147018 363012 147024
rect 363512 4888 363564 4894
rect 363512 4830 363564 4836
rect 362868 4480 362920 4486
rect 362868 4422 362920 4428
rect 362316 4004 362368 4010
rect 362316 3946 362368 3952
rect 361488 3256 361540 3262
rect 361488 3198 361540 3204
rect 362328 480 362356 3946
rect 363524 480 363552 4830
rect 364168 4690 364196 150470
rect 364444 148442 364472 150484
rect 365102 150470 365668 150498
rect 364432 148436 364484 148442
rect 364432 148378 364484 148384
rect 364248 147688 364300 147694
rect 364248 147630 364300 147636
rect 364156 4684 364208 4690
rect 364156 4626 364208 4632
rect 364260 3330 364288 147630
rect 364616 4956 364668 4962
rect 364616 4898 364668 4904
rect 364248 3324 364300 3330
rect 364248 3266 364300 3272
rect 364628 480 364656 4898
rect 365640 4146 365668 150470
rect 365824 147694 365852 150484
rect 366482 150470 366956 150498
rect 366928 147778 366956 150470
rect 366928 147750 367140 147778
rect 365812 147688 365864 147694
rect 365812 147630 365864 147636
rect 367008 147688 367060 147694
rect 367008 147630 367060 147636
rect 367020 6914 367048 147630
rect 367112 147014 367140 147750
rect 367204 147694 367232 150484
rect 367862 150470 368336 150498
rect 367192 147688 367244 147694
rect 367192 147630 367244 147636
rect 367100 147008 367152 147014
rect 367100 146950 367152 146956
rect 366928 6886 367048 6914
rect 366928 4622 366956 6886
rect 368204 5092 368256 5098
rect 368204 5034 368256 5040
rect 367008 5024 367060 5030
rect 367008 4966 367060 4972
rect 366916 4616 366968 4622
rect 366916 4558 366968 4564
rect 365628 4140 365680 4146
rect 365628 4082 365680 4088
rect 365812 3936 365864 3942
rect 365812 3878 365864 3884
rect 365824 480 365852 3878
rect 367020 480 367048 4966
rect 368216 480 368244 5034
rect 368308 4758 368336 150470
rect 368584 148374 368612 150484
rect 369242 150470 369808 150498
rect 368572 148368 368624 148374
rect 368572 148310 368624 148316
rect 368388 147688 368440 147694
rect 368388 147630 368440 147636
rect 368296 4752 368348 4758
rect 368296 4694 368348 4700
rect 368400 3398 368428 147630
rect 369780 4010 369808 150470
rect 369964 147694 369992 150484
rect 370608 148646 370636 150484
rect 370596 148640 370648 148646
rect 370596 148582 370648 148588
rect 371344 147694 371372 150484
rect 372002 150470 372476 150498
rect 369952 147688 370004 147694
rect 369952 147630 370004 147636
rect 371148 147688 371200 147694
rect 371148 147630 371200 147636
rect 371332 147688 371384 147694
rect 371332 147630 371384 147636
rect 370136 15904 370188 15910
rect 370136 15846 370188 15852
rect 369768 4004 369820 4010
rect 369768 3946 369820 3952
rect 369400 3868 369452 3874
rect 369400 3810 369452 3816
rect 368388 3392 368440 3398
rect 368388 3334 368440 3340
rect 369412 480 369440 3810
rect 370148 490 370176 15846
rect 371160 5506 371188 147630
rect 371240 18624 371292 18630
rect 371240 18566 371292 18572
rect 371148 5500 371200 5506
rect 371148 5442 371200 5448
rect 370424 598 370636 626
rect 370424 490 370452 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370148 462 370452 490
rect 370608 480 370636 598
rect 371252 490 371280 18566
rect 372448 5438 372476 150470
rect 372632 149054 372660 150484
rect 373382 150470 373948 150498
rect 372620 149048 372672 149054
rect 372620 148990 372672 148996
rect 372528 147688 372580 147694
rect 372528 147630 372580 147636
rect 372436 5432 372488 5438
rect 372436 5374 372488 5380
rect 372540 4078 372568 147630
rect 372528 4072 372580 4078
rect 372528 4014 372580 4020
rect 373920 3942 373948 150470
rect 374012 147694 374040 150484
rect 374762 150470 375236 150498
rect 374644 149048 374696 149054
rect 374644 148990 374696 148996
rect 374000 147688 374052 147694
rect 374000 147630 374052 147636
rect 374656 146946 374684 148990
rect 374644 146940 374696 146946
rect 374644 146882 374696 146888
rect 375208 11762 375236 150470
rect 375392 147694 375420 150484
rect 376142 150470 376616 150498
rect 375288 147688 375340 147694
rect 375288 147630 375340 147636
rect 375380 147688 375432 147694
rect 375380 147630 375432 147636
rect 375196 11756 375248 11762
rect 375196 11698 375248 11704
rect 375196 6588 375248 6594
rect 375196 6530 375248 6536
rect 374092 4820 374144 4826
rect 374092 4762 374144 4768
rect 373908 3936 373960 3942
rect 373908 3878 373960 3884
rect 372896 3732 372948 3738
rect 372896 3674 372948 3680
rect 371528 598 371740 626
rect 371528 490 371556 598
rect 370566 -960 370678 480
rect 371252 462 371556 490
rect 371712 480 371740 598
rect 372908 480 372936 3674
rect 374104 480 374132 4762
rect 375208 3346 375236 6530
rect 375300 5370 375328 147630
rect 375288 5364 375340 5370
rect 375288 5306 375340 5312
rect 376588 5302 376616 150470
rect 376772 147694 376800 150484
rect 377404 148504 377456 148510
rect 377404 148446 377456 148452
rect 376668 147688 376720 147694
rect 376668 147630 376720 147636
rect 376760 147688 376812 147694
rect 376760 147630 376812 147636
rect 376576 5296 376628 5302
rect 376576 5238 376628 5244
rect 376680 3874 376708 147630
rect 377416 4894 377444 148446
rect 377508 147898 377536 150484
rect 377496 147892 377548 147898
rect 377496 147834 377548 147840
rect 378152 147694 378180 150484
rect 378888 148510 378916 150484
rect 378876 148504 378928 148510
rect 378876 148446 378928 148452
rect 379532 147694 379560 150484
rect 380190 150470 380756 150498
rect 378048 147688 378100 147694
rect 378048 147630 378100 147636
rect 378140 147688 378192 147694
rect 378140 147630 378192 147636
rect 379428 147688 379480 147694
rect 379428 147630 379480 147636
rect 379520 147688 379572 147694
rect 379520 147630 379572 147636
rect 378060 8974 378088 147630
rect 378140 25560 378192 25566
rect 378140 25502 378192 25508
rect 378152 16574 378180 25502
rect 378152 16546 378456 16574
rect 377680 8968 377732 8974
rect 377680 8910 377732 8916
rect 378048 8968 378100 8974
rect 378048 8910 378100 8916
rect 377404 4888 377456 4894
rect 377404 4830 377456 4836
rect 376668 3868 376720 3874
rect 376668 3810 376720 3816
rect 376484 3800 376536 3806
rect 376484 3742 376536 3748
rect 375208 3318 375328 3346
rect 375300 480 375328 3318
rect 376496 480 376524 3742
rect 377692 480 377720 8910
rect 378428 490 378456 16546
rect 379440 5234 379468 147630
rect 379428 5228 379480 5234
rect 379428 5170 379480 5176
rect 380728 5166 380756 150470
rect 380912 147694 380940 150484
rect 381570 150470 382228 150498
rect 380808 147688 380860 147694
rect 380808 147630 380860 147636
rect 380900 147688 380952 147694
rect 380900 147630 380952 147636
rect 382096 147688 382148 147694
rect 382096 147630 382148 147636
rect 380716 5160 380768 5166
rect 380716 5102 380768 5108
rect 380820 3806 380848 147630
rect 382108 7886 382136 147630
rect 382096 7880 382148 7886
rect 382096 7822 382148 7828
rect 381176 6520 381228 6526
rect 381176 6462 381228 6468
rect 380808 3800 380860 3806
rect 380808 3742 380860 3748
rect 379980 3528 380032 3534
rect 379980 3470 380032 3476
rect 378704 598 378916 626
rect 378704 490 378732 598
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 462 378732 490
rect 378888 480 378916 598
rect 379992 480 380020 3470
rect 381188 480 381216 6462
rect 382200 3738 382228 150470
rect 382292 147694 382320 150484
rect 382950 150470 383516 150498
rect 382280 147688 382332 147694
rect 382280 147630 382332 147636
rect 383488 17270 383516 150470
rect 383672 147694 383700 150484
rect 384330 150470 384896 150498
rect 383568 147688 383620 147694
rect 383568 147630 383620 147636
rect 383660 147688 383712 147694
rect 383660 147630 383712 147636
rect 383476 17264 383528 17270
rect 383476 17206 383528 17212
rect 382372 6452 382424 6458
rect 382372 6394 382424 6400
rect 382188 3732 382240 3738
rect 382188 3674 382240 3680
rect 382384 480 382412 6394
rect 383580 5098 383608 147630
rect 383568 5092 383620 5098
rect 383568 5034 383620 5040
rect 384868 4962 384896 150470
rect 385052 147830 385080 150484
rect 385710 150470 386368 150498
rect 385224 148980 385276 148986
rect 385224 148922 385276 148928
rect 385040 147824 385092 147830
rect 385040 147766 385092 147772
rect 384948 147688 385000 147694
rect 384948 147630 385000 147636
rect 384856 4956 384908 4962
rect 384856 4898 384908 4904
rect 384764 4888 384816 4894
rect 384764 4830 384816 4836
rect 383568 3664 383620 3670
rect 383568 3606 383620 3612
rect 383580 480 383608 3606
rect 384776 480 384804 4830
rect 384960 3670 384988 147630
rect 385236 16574 385264 148922
rect 385236 16546 386000 16574
rect 384948 3664 385000 3670
rect 384948 3606 385000 3612
rect 385972 480 386000 16546
rect 386340 3534 386368 150470
rect 386432 147694 386460 150484
rect 387076 148034 387104 150484
rect 387064 148028 387116 148034
rect 387064 147970 387116 147976
rect 387812 147694 387840 150484
rect 388470 150470 389036 150498
rect 388076 148912 388128 148918
rect 388076 148854 388128 148860
rect 386420 147688 386472 147694
rect 386420 147630 386472 147636
rect 387708 147688 387760 147694
rect 387708 147630 387760 147636
rect 387800 147688 387852 147694
rect 387800 147630 387852 147636
rect 387720 5030 387748 147630
rect 388088 16574 388116 148854
rect 388088 16546 388300 16574
rect 387708 5024 387760 5030
rect 387708 4966 387760 4972
rect 386328 3528 386380 3534
rect 386328 3470 386380 3476
rect 387156 3460 387208 3466
rect 387156 3402 387208 3408
rect 387168 480 387196 3402
rect 388272 480 388300 16546
rect 389008 4894 389036 150470
rect 389100 147778 389128 150484
rect 389732 148844 389784 148850
rect 389732 148786 389784 148792
rect 389100 147762 389220 147778
rect 389100 147756 389232 147762
rect 389100 147750 389180 147756
rect 389180 147698 389232 147704
rect 389088 147688 389140 147694
rect 389088 147630 389140 147636
rect 388996 4888 389048 4894
rect 388996 4830 389048 4836
rect 389100 3466 389128 147630
rect 389744 142154 389772 148786
rect 389836 147966 389864 150484
rect 390100 148028 390152 148034
rect 390100 147970 390152 147976
rect 389824 147960 389876 147966
rect 389824 147902 389876 147908
rect 390112 145586 390140 147970
rect 390100 145580 390152 145586
rect 390100 145522 390152 145528
rect 389744 142126 389864 142154
rect 389456 6384 389508 6390
rect 389456 6326 389508 6332
rect 389088 3460 389140 3466
rect 389088 3402 389140 3408
rect 389468 480 389496 6326
rect 389836 4214 389864 142126
rect 390480 4826 390508 150484
rect 391216 147694 391244 150484
rect 391204 147688 391256 147694
rect 391204 147630 391256 147636
rect 391860 6914 391888 150484
rect 392610 150470 393176 150498
rect 392584 147688 392636 147694
rect 392584 147630 392636 147636
rect 392596 7818 392624 147630
rect 393148 142154 393176 150470
rect 393240 145994 393268 150484
rect 393504 148776 393556 148782
rect 393504 148718 393556 148724
rect 393228 145988 393280 145994
rect 393228 145930 393280 145936
rect 393148 142126 393268 142154
rect 392584 7812 392636 7818
rect 392584 7754 392636 7760
rect 391768 6886 391888 6914
rect 390468 4820 390520 4826
rect 390468 4762 390520 4768
rect 389824 4208 389876 4214
rect 389824 4150 389876 4156
rect 391768 3602 391796 6886
rect 393044 6316 393096 6322
rect 393044 6258 393096 6264
rect 391848 4208 391900 4214
rect 391848 4150 391900 4156
rect 390652 3596 390704 3602
rect 390652 3538 390704 3544
rect 391756 3596 391808 3602
rect 391756 3538 391808 3544
rect 390664 480 390692 3538
rect 391860 480 391888 4150
rect 393056 480 393084 6258
rect 393240 5914 393268 142126
rect 393516 16574 393544 148718
rect 393976 148102 394004 150484
rect 393964 148096 394016 148102
rect 393964 148038 394016 148044
rect 393516 16546 394280 16574
rect 393228 5908 393280 5914
rect 393228 5850 393280 5856
rect 394252 480 394280 16546
rect 394620 5982 394648 150484
rect 395370 150470 395936 150498
rect 395908 15910 395936 150470
rect 395896 15904 395948 15910
rect 395896 15846 395948 15852
rect 394608 5976 394660 5982
rect 394608 5918 394660 5924
rect 395344 4276 395396 4282
rect 395344 4218 395396 4224
rect 395356 480 395384 4218
rect 396000 2854 396028 150484
rect 396644 147694 396672 150484
rect 397288 150470 397394 150498
rect 396632 147688 396684 147694
rect 396632 147630 396684 147636
rect 397288 33794 397316 150470
rect 398024 148238 398052 150484
rect 398012 148232 398064 148238
rect 398012 148174 398064 148180
rect 397368 147688 397420 147694
rect 397368 147630 397420 147636
rect 397276 33788 397328 33794
rect 397276 33730 397328 33736
rect 396540 6180 396592 6186
rect 396540 6122 396592 6128
rect 395988 2848 396040 2854
rect 395988 2790 396040 2796
rect 396552 480 396580 6122
rect 397380 6050 397408 147630
rect 398760 6798 398788 150484
rect 399418 150470 400076 150498
rect 400048 7750 400076 150470
rect 400036 7744 400088 7750
rect 400036 7686 400088 7692
rect 398748 6792 398800 6798
rect 398748 6734 398800 6740
rect 400036 6248 400088 6254
rect 400036 6190 400088 6196
rect 397368 6044 397420 6050
rect 397368 5986 397420 5992
rect 398932 4412 398984 4418
rect 398932 4354 398984 4360
rect 397736 3120 397788 3126
rect 397736 3062 397788 3068
rect 397748 480 397776 3062
rect 398944 480 398972 4354
rect 400048 2802 400076 6190
rect 400140 2922 400168 150484
rect 400404 148708 400456 148714
rect 400404 148650 400456 148656
rect 400416 16574 400444 148650
rect 400784 147694 400812 150484
rect 401520 148034 401548 150484
rect 402164 148306 402192 150484
rect 402152 148300 402204 148306
rect 402152 148242 402204 148248
rect 402900 148170 402928 150484
rect 402888 148164 402940 148170
rect 402888 148106 402940 148112
rect 401508 148028 401560 148034
rect 401508 147970 401560 147976
rect 403544 147694 403572 150484
rect 404188 150470 404294 150498
rect 400772 147688 400824 147694
rect 400772 147630 400824 147636
rect 401508 147688 401560 147694
rect 401508 147630 401560 147636
rect 403532 147688 403584 147694
rect 403532 147630 403584 147636
rect 400416 16546 400904 16574
rect 400128 2916 400180 2922
rect 400128 2858 400180 2864
rect 400048 2774 400168 2802
rect 400140 480 400168 2774
rect 400876 490 400904 16546
rect 401520 6118 401548 147630
rect 404188 145926 404216 150470
rect 404924 147694 404952 150484
rect 405582 150470 405688 150498
rect 404268 147688 404320 147694
rect 404268 147630 404320 147636
rect 404912 147688 404964 147694
rect 404912 147630 404964 147636
rect 404176 145920 404228 145926
rect 404176 145862 404228 145868
rect 403624 7608 403676 7614
rect 403624 7550 403676 7556
rect 401508 6112 401560 6118
rect 401508 6054 401560 6060
rect 402520 4344 402572 4350
rect 402520 4286 402572 4292
rect 401152 598 401364 626
rect 401152 490 401180 598
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 462 401180 490
rect 401336 480 401364 598
rect 402532 480 402560 4286
rect 403636 480 403664 7550
rect 404280 6730 404308 147630
rect 404268 6724 404320 6730
rect 404268 6666 404320 6672
rect 405660 6662 405688 150470
rect 406304 149054 406332 150484
rect 406962 150470 407068 150498
rect 407698 150470 408264 150498
rect 406292 149048 406344 149054
rect 406292 148990 406344 148996
rect 406384 148572 406436 148578
rect 406384 148514 406436 148520
rect 405648 6656 405700 6662
rect 405648 6598 405700 6604
rect 406396 5574 406424 148514
rect 407040 7682 407068 150470
rect 408236 142154 408264 150470
rect 408328 144226 408356 150484
rect 409064 148714 409092 150484
rect 409722 150470 409828 150498
rect 409052 148708 409104 148714
rect 409052 148650 409104 148656
rect 408316 144220 408368 144226
rect 408316 144162 408368 144168
rect 408236 142126 408448 142154
rect 407028 7676 407080 7682
rect 407028 7618 407080 7624
rect 408420 6594 408448 142126
rect 408408 6588 408460 6594
rect 408408 6530 408460 6536
rect 409800 6526 409828 150470
rect 410444 148986 410472 150484
rect 411102 150470 411208 150498
rect 410432 148980 410484 148986
rect 410432 148922 410484 148928
rect 410800 148708 410852 148714
rect 410800 148650 410852 148656
rect 410812 147558 410840 148650
rect 410800 147552 410852 147558
rect 410800 147494 410852 147500
rect 409880 147076 409932 147082
rect 409880 147018 409932 147024
rect 409892 16574 409920 147018
rect 409892 16546 410840 16574
rect 409788 6520 409840 6526
rect 409788 6462 409840 6468
rect 406384 5568 406436 5574
rect 406384 5510 406436 5516
rect 407212 5568 407264 5574
rect 407212 5510 407264 5516
rect 406016 4548 406068 4554
rect 406016 4490 406068 4496
rect 404820 3188 404872 3194
rect 404820 3130 404872 3136
rect 404832 480 404860 3130
rect 406028 480 406056 4490
rect 407224 480 407252 5510
rect 409604 4480 409656 4486
rect 409604 4422 409656 4428
rect 408408 3256 408460 3262
rect 408408 3198 408460 3204
rect 408420 480 408448 3198
rect 409616 480 409644 4422
rect 410812 480 410840 16546
rect 411180 7614 411208 150470
rect 411824 147694 411852 150484
rect 411812 147688 411864 147694
rect 411812 147630 411864 147636
rect 412468 18630 412496 150484
rect 413112 148850 413140 150484
rect 413862 150470 413968 150498
rect 413100 148844 413152 148850
rect 413100 148786 413152 148792
rect 413284 148436 413336 148442
rect 413284 148378 413336 148384
rect 412548 147688 412600 147694
rect 412548 147630 412600 147636
rect 412456 18624 412508 18630
rect 412456 18566 412508 18572
rect 411168 7608 411220 7614
rect 411168 7550 411220 7556
rect 412560 6458 412588 147630
rect 413296 13734 413324 148378
rect 413284 13728 413336 13734
rect 413284 13670 413336 13676
rect 412548 6452 412600 6458
rect 412548 6394 412600 6400
rect 413940 6390 413968 150470
rect 414492 148782 414520 150484
rect 415242 150470 415348 150498
rect 414480 148776 414532 148782
rect 414480 148718 414532 148724
rect 414664 148640 414716 148646
rect 414664 148582 414716 148588
rect 414296 13728 414348 13734
rect 414296 13670 414348 13676
rect 413928 6384 413980 6390
rect 413928 6326 413980 6332
rect 413100 4684 413152 4690
rect 413100 4626 413152 4632
rect 411904 3324 411956 3330
rect 411904 3266 411956 3272
rect 411916 480 411944 3266
rect 413112 480 413140 4626
rect 414308 480 414336 13670
rect 414676 7954 414704 148582
rect 415320 13122 415348 150470
rect 415872 147694 415900 150484
rect 416622 150470 416728 150498
rect 415860 147688 415912 147694
rect 415860 147630 415912 147636
rect 416596 147688 416648 147694
rect 416596 147630 416648 147636
rect 415308 13116 415360 13122
rect 415308 13058 415360 13064
rect 414664 7948 414716 7954
rect 414664 7890 414716 7896
rect 416608 6322 416636 147630
rect 416700 147490 416728 150470
rect 417252 148714 417280 150484
rect 418002 150470 418108 150498
rect 417240 148708 417292 148714
rect 417240 148650 417292 148656
rect 416688 147484 416740 147490
rect 416688 147426 416740 147432
rect 416780 147008 416832 147014
rect 416780 146950 416832 146956
rect 416792 16574 416820 146950
rect 416792 16546 417464 16574
rect 416596 6316 416648 6322
rect 416596 6258 416648 6264
rect 416688 4616 416740 4622
rect 416688 4558 416740 4564
rect 415492 4140 415544 4146
rect 415492 4082 415544 4088
rect 415504 480 415532 4082
rect 416700 480 416728 4558
rect 417436 490 417464 16546
rect 418080 6254 418108 150470
rect 418632 148646 418660 150484
rect 419382 150470 419488 150498
rect 418620 148640 418672 148646
rect 418620 148582 418672 148588
rect 418804 148368 418856 148374
rect 418804 148310 418856 148316
rect 418068 6248 418120 6254
rect 418068 6190 418120 6196
rect 418816 4214 418844 148310
rect 419460 10334 419488 150470
rect 420012 148918 420040 150484
rect 420762 150470 420868 150498
rect 420000 148912 420052 148918
rect 420000 148854 420052 148860
rect 419448 10328 419500 10334
rect 419448 10270 419500 10276
rect 420184 4752 420236 4758
rect 420184 4694 420236 4700
rect 418804 4208 418856 4214
rect 418804 4150 418856 4156
rect 418988 3392 419040 3398
rect 418988 3334 419040 3340
rect 417712 598 417924 626
rect 417712 490 417740 598
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 462 417740 490
rect 417896 480 417924 598
rect 419000 480 419028 3334
rect 420196 480 420224 4694
rect 420840 2990 420868 150470
rect 421392 147694 421420 150484
rect 422050 150470 422156 150498
rect 421380 147688 421432 147694
rect 421380 147630 421432 147636
rect 422128 6186 422156 150470
rect 422772 148578 422800 150484
rect 423430 150470 423628 150498
rect 422760 148572 422812 148578
rect 422760 148514 422812 148520
rect 422208 147688 422260 147694
rect 422208 147630 422260 147636
rect 422116 6180 422168 6186
rect 422116 6122 422168 6128
rect 422220 4282 422248 147630
rect 423600 4350 423628 150470
rect 424152 147694 424180 150484
rect 424810 150470 425008 150498
rect 425546 150470 426020 150498
rect 424140 147688 424192 147694
rect 424140 147630 424192 147636
rect 424876 7948 424928 7954
rect 424876 7890 424928 7896
rect 423772 5500 423824 5506
rect 423772 5442 423824 5448
rect 423588 4344 423640 4350
rect 423588 4286 423640 4292
rect 422208 4276 422260 4282
rect 422208 4218 422260 4224
rect 421380 4208 421432 4214
rect 421380 4150 421432 4156
rect 420828 2984 420880 2990
rect 420828 2926 420880 2932
rect 421392 480 421420 4150
rect 422576 4004 422628 4010
rect 422576 3946 422628 3952
rect 422588 480 422616 3946
rect 423784 480 423812 5442
rect 424784 4140 424836 4146
rect 424784 4082 424836 4088
rect 424796 3058 424824 4082
rect 424888 3482 424916 7890
rect 424980 4146 425008 150470
rect 425704 148504 425756 148510
rect 425704 148446 425756 148452
rect 425716 8022 425744 148446
rect 425992 142154 426020 150470
rect 426176 147422 426204 150484
rect 426912 147694 426940 150484
rect 427570 150470 427676 150498
rect 426900 147688 426952 147694
rect 426900 147630 426952 147636
rect 426164 147416 426216 147422
rect 426164 147358 426216 147364
rect 425992 142126 426296 142154
rect 425704 8016 425756 8022
rect 425704 7958 425756 7964
rect 426268 4418 426296 142126
rect 427268 5432 427320 5438
rect 427268 5374 427320 5380
rect 426256 4412 426308 4418
rect 426256 4354 426308 4360
rect 424968 4140 425020 4146
rect 424968 4082 425020 4088
rect 426164 4072 426216 4078
rect 426164 4014 426216 4020
rect 424888 3454 425008 3482
rect 424784 3052 424836 3058
rect 424784 2994 424836 3000
rect 424980 480 425008 3454
rect 426176 480 426204 4014
rect 427280 480 427308 5374
rect 427648 4554 427676 150470
rect 428292 148510 428320 150484
rect 428950 150470 429148 150498
rect 428280 148504 428332 148510
rect 428280 148446 428332 148452
rect 427728 147688 427780 147694
rect 427728 147630 427780 147636
rect 427636 4548 427688 4554
rect 427636 4490 427688 4496
rect 427740 3126 427768 147630
rect 427820 146940 427872 146946
rect 427820 146882 427872 146888
rect 427832 16574 427860 146882
rect 427832 16546 428504 16574
rect 427728 3120 427780 3126
rect 427728 3062 427780 3068
rect 428476 480 428504 16546
rect 429120 3194 429148 150470
rect 429580 147694 429608 150484
rect 430316 148442 430344 150484
rect 430304 148436 430356 148442
rect 430304 148378 430356 148384
rect 429844 147824 429896 147830
rect 429844 147766 429896 147772
rect 429568 147688 429620 147694
rect 429568 147630 429620 147636
rect 429856 14482 429884 147766
rect 430960 147762 430988 150484
rect 431710 150470 431816 150498
rect 432354 150470 432736 150498
rect 433090 150470 433288 150498
rect 430948 147756 431000 147762
rect 430948 147698 431000 147704
rect 430488 147688 430540 147694
rect 430488 147630 430540 147636
rect 429844 14476 429896 14482
rect 429844 14418 429896 14424
rect 430500 4486 430528 147630
rect 430856 5364 430908 5370
rect 430856 5306 430908 5312
rect 430488 4480 430540 4486
rect 430488 4422 430540 4428
rect 429660 3936 429712 3942
rect 429660 3878 429712 3884
rect 429108 3188 429160 3194
rect 429108 3130 429160 3136
rect 429672 480 429700 3878
rect 430868 480 430896 5306
rect 431788 4690 431816 150470
rect 432708 148374 432736 150470
rect 432604 148368 432656 148374
rect 432604 148310 432656 148316
rect 432696 148368 432748 148374
rect 432696 148310 432748 148316
rect 431868 147756 431920 147762
rect 431868 147698 431920 147704
rect 431776 4684 431828 4690
rect 431776 4626 431828 4632
rect 431880 3262 431908 147698
rect 432052 11756 432104 11762
rect 432052 11698 432104 11704
rect 431868 3256 431920 3262
rect 431868 3198 431920 3204
rect 432064 480 432092 11698
rect 432616 7954 432644 148310
rect 432604 7948 432656 7954
rect 432604 7890 432656 7896
rect 433260 6914 433288 150470
rect 433720 147762 433748 150484
rect 434456 147830 434484 150484
rect 434444 147824 434496 147830
rect 434444 147766 434496 147772
rect 435100 147762 435128 150484
rect 435850 150470 435956 150498
rect 433708 147756 433760 147762
rect 433708 147698 433760 147704
rect 434628 147756 434680 147762
rect 434628 147698 434680 147704
rect 435088 147756 435140 147762
rect 435088 147698 435140 147704
rect 433168 6886 433288 6914
rect 433168 3330 433196 6886
rect 434444 5296 434496 5302
rect 434444 5238 434496 5244
rect 433248 3868 433300 3874
rect 433248 3810 433300 3816
rect 433156 3324 433208 3330
rect 433156 3266 433208 3272
rect 433260 480 433288 3810
rect 434456 480 434484 5238
rect 434640 4622 434668 147698
rect 435548 8968 435600 8974
rect 435548 8910 435600 8916
rect 434628 4616 434680 4622
rect 434628 4558 434680 4564
rect 435560 480 435588 8910
rect 435928 5506 435956 150470
rect 436100 147892 436152 147898
rect 436100 147834 436152 147840
rect 436008 147756 436060 147762
rect 436008 147698 436060 147704
rect 435916 5500 435968 5506
rect 435916 5442 435968 5448
rect 436020 3398 436048 147698
rect 436112 16574 436140 147834
rect 436480 147354 436508 150484
rect 437230 150470 437336 150498
rect 436468 147348 436520 147354
rect 436468 147290 436520 147296
rect 436112 16546 436784 16574
rect 436008 3392 436060 3398
rect 436008 3334 436060 3340
rect 436756 480 436784 16546
rect 437308 4146 437336 150470
rect 437860 147762 437888 150484
rect 437848 147756 437900 147762
rect 437848 147698 437900 147704
rect 438504 147286 438532 150484
rect 439240 147762 439268 150484
rect 439898 150470 440096 150498
rect 438676 147756 438728 147762
rect 438676 147698 438728 147704
rect 439228 147756 439280 147762
rect 439228 147698 439280 147704
rect 438492 147280 438544 147286
rect 438492 147222 438544 147228
rect 437940 5228 437992 5234
rect 437940 5170 437992 5176
rect 437296 4140 437348 4146
rect 437296 4082 437348 4088
rect 437952 480 437980 5170
rect 438688 4758 438716 147698
rect 439136 8016 439188 8022
rect 439136 7958 439188 7964
rect 438676 4752 438728 4758
rect 438676 4694 438728 4700
rect 439148 480 439176 7958
rect 440068 5438 440096 150470
rect 440148 147756 440200 147762
rect 440148 147698 440200 147704
rect 440056 5432 440108 5438
rect 440056 5374 440108 5380
rect 440160 4078 440188 147698
rect 440620 147218 440648 150484
rect 441278 150470 441476 150498
rect 440608 147212 440660 147218
rect 440608 147154 440660 147160
rect 440148 4072 440200 4078
rect 440148 4014 440200 4020
rect 441448 4010 441476 150470
rect 442000 147762 442028 150484
rect 441988 147756 442040 147762
rect 441988 147698 442040 147704
rect 442644 147150 442672 150484
rect 443380 147762 443408 150484
rect 444038 150470 444236 150498
rect 442816 147756 442868 147762
rect 442816 147698 442868 147704
rect 443368 147756 443420 147762
rect 443368 147698 443420 147704
rect 442632 147144 442684 147150
rect 442632 147086 442684 147092
rect 442632 7880 442684 7886
rect 442632 7822 442684 7828
rect 441528 5160 441580 5166
rect 441528 5102 441580 5108
rect 441436 4004 441488 4010
rect 441436 3946 441488 3952
rect 440332 3800 440384 3806
rect 440332 3742 440384 3748
rect 440344 480 440372 3742
rect 441540 480 441568 5102
rect 442644 480 442672 7822
rect 442828 5370 442856 147698
rect 442816 5364 442868 5370
rect 442816 5306 442868 5312
rect 444208 5302 444236 150470
rect 444288 147756 444340 147762
rect 444288 147698 444340 147704
rect 444196 5296 444248 5302
rect 444196 5238 444248 5244
rect 444300 3942 444328 147698
rect 444760 147082 444788 150484
rect 445418 150470 445616 150498
rect 444748 147076 444800 147082
rect 444748 147018 444800 147024
rect 445024 5092 445076 5098
rect 445024 5034 445076 5040
rect 444288 3936 444340 3942
rect 444288 3878 444340 3884
rect 443828 3732 443880 3738
rect 443828 3674 443880 3680
rect 443840 480 443868 3674
rect 445036 480 445064 5034
rect 445588 3874 445616 150470
rect 446048 147762 446076 150484
rect 446036 147756 446088 147762
rect 446036 147698 446088 147704
rect 446784 145790 446812 150484
rect 447428 147762 447456 150484
rect 448178 150470 448376 150498
rect 447048 147756 447100 147762
rect 447048 147698 447100 147704
rect 447416 147756 447468 147762
rect 447416 147698 447468 147704
rect 446772 145784 446824 145790
rect 446772 145726 446824 145732
rect 445760 17264 445812 17270
rect 445760 17206 445812 17212
rect 445576 3868 445628 3874
rect 445576 3810 445628 3816
rect 445772 490 445800 17206
rect 447060 5234 447088 147698
rect 447048 5228 447100 5234
rect 447048 5170 447100 5176
rect 448348 5166 448376 150470
rect 448428 147756 448480 147762
rect 448428 147698 448480 147704
rect 448336 5160 448388 5166
rect 448336 5102 448388 5108
rect 448440 3806 448468 147698
rect 448808 145858 448836 150484
rect 449558 150470 449848 150498
rect 448796 145852 448848 145858
rect 448796 145794 448848 145800
rect 448520 14476 448572 14482
rect 448520 14418 448572 14424
rect 448428 3800 448480 3806
rect 448428 3742 448480 3748
rect 447416 3664 447468 3670
rect 447416 3606 447468 3612
rect 446048 598 446260 626
rect 446048 490 446076 598
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 462 446076 490
rect 446232 480 446260 598
rect 447428 480 447456 3606
rect 448532 2786 448560 14418
rect 449820 6914 449848 150470
rect 450188 147762 450216 150484
rect 450176 147756 450228 147762
rect 450176 147698 450228 147704
rect 450924 145722 450952 150484
rect 451568 147762 451596 150484
rect 452318 150470 452516 150498
rect 451188 147756 451240 147762
rect 451188 147698 451240 147704
rect 451556 147756 451608 147762
rect 451556 147698 451608 147704
rect 450912 145716 450964 145722
rect 450912 145658 450964 145664
rect 449728 6886 449848 6914
rect 448612 4956 448664 4962
rect 448612 4898 448664 4904
rect 448520 2780 448572 2786
rect 448520 2722 448572 2728
rect 448624 480 448652 4898
rect 449728 3738 449756 6886
rect 451200 5098 451228 147698
rect 451188 5092 451240 5098
rect 451188 5034 451240 5040
rect 452488 5030 452516 150470
rect 452568 147756 452620 147762
rect 452568 147698 452620 147704
rect 452108 5024 452160 5030
rect 452108 4966 452160 4972
rect 452476 5024 452528 5030
rect 452476 4966 452528 4972
rect 449716 3732 449768 3738
rect 449716 3674 449768 3680
rect 450912 3528 450964 3534
rect 450912 3470 450964 3476
rect 449808 2780 449860 2786
rect 449808 2722 449860 2728
rect 449820 480 449848 2722
rect 450924 480 450952 3470
rect 452120 480 452148 4966
rect 452580 3670 452608 147698
rect 452948 145654 452976 150484
rect 453698 150470 453988 150498
rect 452936 145648 452988 145654
rect 452936 145590 452988 145596
rect 452660 145580 452712 145586
rect 452660 145522 452712 145528
rect 452672 16574 452700 145522
rect 452672 16546 453344 16574
rect 452568 3664 452620 3670
rect 452568 3606 452620 3612
rect 453316 480 453344 16546
rect 453960 3534 453988 150470
rect 454328 147762 454356 150484
rect 454316 147756 454368 147762
rect 454316 147698 454368 147704
rect 454972 147014 455000 150484
rect 455708 147762 455736 150484
rect 456366 150470 456656 150498
rect 455236 147756 455288 147762
rect 455236 147698 455288 147704
rect 455696 147756 455748 147762
rect 455696 147698 455748 147704
rect 454960 147008 455012 147014
rect 454960 146950 455012 146956
rect 455248 4962 455276 147698
rect 455236 4956 455288 4962
rect 455236 4898 455288 4904
rect 456628 4826 456656 150470
rect 456800 147960 456852 147966
rect 456800 147902 456852 147908
rect 456708 147756 456760 147762
rect 456708 147698 456760 147704
rect 455696 4820 455748 4826
rect 455696 4762 455748 4768
rect 456616 4820 456668 4826
rect 456616 4762 456668 4768
rect 453948 3528 454000 3534
rect 453948 3470 454000 3476
rect 454500 3460 454552 3466
rect 454500 3402 454552 3408
rect 454512 480 454540 3402
rect 455708 480 455736 4762
rect 456616 3528 456668 3534
rect 456614 3496 456616 3505
rect 456668 3496 456670 3505
rect 456720 3466 456748 147698
rect 456812 3534 456840 147902
rect 457088 146946 457116 150484
rect 457746 150470 458036 150498
rect 457076 146940 457128 146946
rect 457076 146882 457128 146888
rect 456892 7948 456944 7954
rect 456892 7890 456944 7896
rect 456800 3528 456852 3534
rect 456800 3470 456852 3476
rect 456614 3431 456670 3440
rect 456708 3460 456760 3466
rect 456708 3402 456760 3408
rect 456904 480 456932 7890
rect 458008 3777 458036 150470
rect 458468 147762 458496 150484
rect 458456 147756 458508 147762
rect 458456 147698 458508 147704
rect 459112 145586 459140 150484
rect 459848 147762 459876 150484
rect 460506 150470 460796 150498
rect 459468 147756 459520 147762
rect 459468 147698 459520 147704
rect 459836 147756 459888 147762
rect 459836 147698 459888 147704
rect 459100 145580 459152 145586
rect 459100 145522 459152 145528
rect 459480 4894 459508 147698
rect 460388 7812 460440 7818
rect 460388 7754 460440 7760
rect 459192 4888 459244 4894
rect 459192 4830 459244 4836
rect 459468 4888 459520 4894
rect 459468 4830 459520 4836
rect 457994 3768 458050 3777
rect 457994 3703 458050 3712
rect 458088 3528 458140 3534
rect 458180 3528 458232 3534
rect 458088 3470 458140 3476
rect 458178 3496 458180 3505
rect 458232 3496 458234 3505
rect 458100 480 458128 3470
rect 458178 3431 458234 3440
rect 459204 480 459232 4830
rect 460400 480 460428 7754
rect 460768 3505 460796 150470
rect 460848 147756 460900 147762
rect 460848 147698 460900 147704
rect 460860 3641 460888 147698
rect 461228 147694 461256 150484
rect 461886 150470 462176 150498
rect 461216 147688 461268 147694
rect 461216 147630 461268 147636
rect 460846 3632 460902 3641
rect 460846 3567 460902 3576
rect 461584 3596 461636 3602
rect 461584 3538 461636 3544
rect 460754 3496 460810 3505
rect 460754 3431 460810 3440
rect 461596 480 461624 3538
rect 462148 3369 462176 150470
rect 465080 148096 465132 148102
rect 465080 148038 465132 148044
rect 464344 147756 464396 147762
rect 464344 147698 464396 147704
rect 462228 147688 462280 147694
rect 462228 147630 462280 147636
rect 462240 3602 462268 147630
rect 463700 145988 463752 145994
rect 463700 145930 463752 145936
rect 463712 16574 463740 145930
rect 463712 16546 464016 16574
rect 462780 5908 462832 5914
rect 462780 5850 462832 5856
rect 462228 3596 462280 3602
rect 462228 3538 462280 3544
rect 462134 3360 462190 3369
rect 462134 3295 462190 3304
rect 462792 480 462820 5850
rect 463988 480 464016 16546
rect 464356 7886 464384 147698
rect 465092 16574 465120 148038
rect 468484 148028 468536 148034
rect 468484 147970 468536 147976
rect 467104 147824 467156 147830
rect 467104 147766 467156 147772
rect 465092 16546 465212 16574
rect 464344 7880 464396 7886
rect 464344 7822 464396 7828
rect 465184 480 465212 16546
rect 467116 7818 467144 147766
rect 467472 15904 467524 15910
rect 467472 15846 467524 15852
rect 467104 7812 467156 7818
rect 467104 7754 467156 7760
rect 466276 5976 466328 5982
rect 466276 5918 466328 5924
rect 466288 480 466316 5918
rect 467484 480 467512 15846
rect 468496 7954 468524 147970
rect 470600 33788 470652 33794
rect 470600 33730 470652 33736
rect 468484 7948 468536 7954
rect 468484 7890 468536 7896
rect 469864 6044 469916 6050
rect 469864 5986 469916 5992
rect 468668 2848 468720 2854
rect 468668 2790 468720 2796
rect 468680 480 468708 2790
rect 469876 480 469904 5986
rect 470612 490 470640 33730
rect 471256 33114 471284 557602
rect 472636 153202 472664 559098
rect 475396 179382 475424 560594
rect 479536 219434 479564 560662
rect 482296 259418 482324 560730
rect 483676 313274 483704 560798
rect 485056 365702 485084 560866
rect 486436 419490 486464 561002
rect 558932 560998 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683262 580212 683839
rect 580172 683256 580224 683262
rect 580172 683198 580224 683204
rect 580172 670812 580224 670818
rect 580172 670754 580224 670760
rect 580184 670721 580212 670754
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 558920 560992 558972 560998
rect 558920 560934 558972 560940
rect 497464 559360 497516 559366
rect 497464 559302 497516 559308
rect 490564 559224 490616 559230
rect 490564 559166 490616 559172
rect 489184 557728 489236 557734
rect 489184 557670 489236 557676
rect 486424 419484 486476 419490
rect 486424 419426 486476 419432
rect 485044 365696 485096 365702
rect 485044 365638 485096 365644
rect 483664 313268 483716 313274
rect 483664 313210 483716 313216
rect 482284 259412 482336 259418
rect 482284 259354 482336 259360
rect 479524 219428 479576 219434
rect 479524 219370 479576 219376
rect 489196 193186 489224 557670
rect 490576 233238 490604 559166
rect 493324 557796 493376 557802
rect 493324 557738 493376 557744
rect 493336 273222 493364 557738
rect 497476 325650 497504 559302
rect 522304 559020 522356 559026
rect 522304 558962 522356 558968
rect 500224 558000 500276 558006
rect 500224 557942 500276 557948
rect 500236 379506 500264 557942
rect 500224 379500 500276 379506
rect 500224 379442 500276 379448
rect 497464 325644 497516 325650
rect 497464 325586 497516 325592
rect 493324 273216 493376 273222
rect 493324 273158 493376 273164
rect 490564 233232 490616 233238
rect 490564 233174 490616 233180
rect 522316 206990 522344 558962
rect 580724 557388 580776 557394
rect 580724 557330 580776 557336
rect 580632 557184 580684 557190
rect 580632 557126 580684 557132
rect 580448 557116 580500 557122
rect 580448 557058 580500 557064
rect 580356 556708 580408 556714
rect 580356 556650 580408 556656
rect 580264 556232 580316 556238
rect 580264 556174 580316 556180
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 579620 405680 579672 405686
rect 579620 405622 579672 405628
rect 579632 404977 579660 405622
rect 579618 404968 579674 404977
rect 579618 404903 579674 404912
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 579896 325644 579948 325650
rect 579896 325586 579948 325592
rect 579908 325281 579936 325586
rect 579894 325272 579950 325281
rect 579894 325207 579950 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 579620 299464 579672 299470
rect 579620 299406 579672 299412
rect 579632 298761 579660 299406
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 579896 219428 579948 219434
rect 579896 219370 579948 219376
rect 579908 219065 579936 219370
rect 579894 219056 579950 219065
rect 579894 218991 579950 219000
rect 522304 206984 522356 206990
rect 522304 206926 522356 206932
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 489184 193180 489236 193186
rect 489184 193122 489236 193128
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 475384 179376 475436 179382
rect 475384 179318 475436 179324
rect 579988 179376 580040 179382
rect 579988 179318 580040 179324
rect 580000 179217 580028 179318
rect 579986 179208 580042 179217
rect 579986 179143 580042 179152
rect 580276 165889 580304 556174
rect 580368 431633 580396 556650
rect 580460 471481 580488 557058
rect 580540 556980 580592 556986
rect 580540 556922 580592 556928
rect 580552 484673 580580 556922
rect 580644 511329 580672 557126
rect 580736 524521 580764 557330
rect 580816 557320 580868 557326
rect 580816 557262 580868 557268
rect 580828 537849 580856 557262
rect 580814 537840 580870 537849
rect 580814 537775 580870 537784
rect 580722 524512 580778 524521
rect 580722 524447 580778 524456
rect 580630 511320 580686 511329
rect 580630 511255 580686 511264
rect 580538 484664 580594 484673
rect 580538 484599 580594 484608
rect 580446 471472 580502 471481
rect 580446 471407 580502 471416
rect 580354 431624 580410 431633
rect 580354 431559 580410 431568
rect 580262 165880 580318 165889
rect 580262 165815 580318 165824
rect 472624 153196 472676 153202
rect 472624 153138 472676 153144
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 485780 149048 485832 149054
rect 485780 148990 485832 148996
rect 478880 148300 478932 148306
rect 478880 148242 478932 148248
rect 471980 148232 472032 148238
rect 471980 148174 472032 148180
rect 471244 33108 471296 33114
rect 471244 33050 471296 33056
rect 471992 16574 472020 148174
rect 475384 148164 475436 148170
rect 475384 148106 475436 148112
rect 471992 16546 472296 16574
rect 470888 598 471100 626
rect 470888 490 470916 598
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 462 470916 490
rect 471072 480 471100 598
rect 472268 480 472296 16546
rect 474556 7744 474608 7750
rect 474556 7686 474608 7692
rect 473452 6792 473504 6798
rect 473452 6734 473504 6740
rect 473464 480 473492 6734
rect 474568 480 474596 7686
rect 475396 5574 475424 148106
rect 478144 7948 478196 7954
rect 478144 7890 478196 7896
rect 476948 6112 477000 6118
rect 476948 6054 477000 6060
rect 475384 5568 475436 5574
rect 475384 5510 475436 5516
rect 475752 2916 475804 2922
rect 475752 2858 475804 2864
rect 475764 480 475792 2858
rect 476960 480 476988 6054
rect 478156 480 478184 7890
rect 478892 490 478920 148242
rect 483020 147620 483072 147626
rect 483020 147562 483072 147568
rect 481640 145920 481692 145926
rect 481640 145862 481692 145868
rect 481652 16574 481680 145862
rect 483032 16574 483060 147562
rect 485792 16574 485820 148990
rect 492680 148980 492732 148986
rect 492680 148922 492732 148928
rect 490012 147552 490064 147558
rect 490012 147494 490064 147500
rect 489184 144220 489236 144226
rect 489184 144162 489236 144168
rect 481652 16546 482416 16574
rect 483032 16546 484072 16574
rect 485792 16546 486464 16574
rect 481732 6724 481784 6730
rect 481732 6666 481784 6672
rect 480536 5568 480588 5574
rect 480536 5510 480588 5516
rect 479168 598 479380 626
rect 479168 490 479196 598
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 478892 462 479196 490
rect 479352 480 479380 598
rect 480548 480 480576 5510
rect 481744 480 481772 6666
rect 482388 490 482416 16546
rect 482664 598 482876 626
rect 482664 490 482692 598
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 462 482692 490
rect 482848 480 482876 598
rect 484044 480 484072 16546
rect 485228 6656 485280 6662
rect 485228 6598 485280 6604
rect 485240 480 485268 6598
rect 486436 480 486464 16546
rect 487620 7676 487672 7682
rect 487620 7618 487672 7624
rect 487632 480 487660 7618
rect 488816 6588 488868 6594
rect 488816 6530 488868 6536
rect 488828 480 488856 6530
rect 489196 2922 489224 144162
rect 490024 16574 490052 147494
rect 492692 16574 492720 148922
rect 504364 148912 504416 148918
rect 504364 148854 504416 148860
rect 497464 148844 497516 148850
rect 497464 148786 497516 148792
rect 496820 18624 496872 18630
rect 496820 18566 496872 18572
rect 496832 16574 496860 18566
rect 490024 16546 490696 16574
rect 492692 16546 493088 16574
rect 496832 16546 497136 16574
rect 489184 2916 489236 2922
rect 489184 2858 489236 2864
rect 489920 2916 489972 2922
rect 489920 2858 489972 2864
rect 489932 480 489960 2858
rect 490668 490 490696 16546
rect 492312 6520 492364 6526
rect 492312 6462 492364 6468
rect 490944 598 491156 626
rect 490944 490 490972 598
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 462 490972 490
rect 491128 480 491156 598
rect 492324 480 492352 6462
rect 493060 490 493088 16546
rect 494704 7608 494756 7614
rect 494704 7550 494756 7556
rect 493336 598 493548 626
rect 493336 490 493364 598
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 462 493364 490
rect 493520 480 493548 598
rect 494716 480 494744 7550
rect 495900 6452 495952 6458
rect 495900 6394 495952 6400
rect 495912 480 495940 6394
rect 497108 480 497136 16546
rect 497476 5574 497504 148786
rect 499580 148776 499632 148782
rect 499580 148718 499632 148724
rect 499592 16574 499620 148718
rect 502984 148708 503036 148714
rect 502984 148650 503036 148656
rect 501604 147484 501656 147490
rect 501604 147426 501656 147432
rect 499592 16546 500632 16574
rect 499396 6384 499448 6390
rect 499396 6326 499448 6332
rect 497464 5568 497516 5574
rect 497464 5510 497516 5516
rect 498200 5568 498252 5574
rect 498200 5510 498252 5516
rect 498212 480 498240 5510
rect 499408 480 499436 6326
rect 500604 480 500632 16546
rect 501328 13116 501380 13122
rect 501328 13058 501380 13064
rect 501340 490 501368 13058
rect 501616 2922 501644 147426
rect 502892 6316 502944 6322
rect 502892 6258 502944 6264
rect 501604 2916 501656 2922
rect 501604 2858 501656 2864
rect 502904 1442 502932 6258
rect 502996 5574 503024 148650
rect 504376 5642 504404 148854
rect 506480 148640 506532 148646
rect 506480 148582 506532 148588
rect 506492 16574 506520 148582
rect 514760 148572 514812 148578
rect 514760 148514 514812 148520
rect 506492 16546 507256 16574
rect 506480 6248 506532 6254
rect 506480 6190 506532 6196
rect 504364 5636 504416 5642
rect 504364 5578 504416 5584
rect 502984 5568 503036 5574
rect 502984 5510 503036 5516
rect 505376 5568 505428 5574
rect 505376 5510 505428 5516
rect 504180 2916 504232 2922
rect 504180 2858 504232 2864
rect 502904 1414 503024 1442
rect 501616 598 501828 626
rect 501616 490 501644 598
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 462 501644 490
rect 501800 480 501828 598
rect 502996 480 503024 1414
rect 504192 480 504220 2858
rect 505388 480 505416 5510
rect 506492 480 506520 6190
rect 507228 490 507256 16546
rect 508872 10328 508924 10334
rect 508872 10270 508924 10276
rect 507504 598 507716 626
rect 507504 490 507532 598
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 462 507532 490
rect 507688 480 507716 598
rect 508884 480 508912 10270
rect 513564 6180 513616 6186
rect 513564 6122 513616 6128
rect 510068 5636 510120 5642
rect 510068 5578 510120 5584
rect 510080 480 510108 5578
rect 512460 4276 512512 4282
rect 512460 4218 512512 4224
rect 511264 2984 511316 2990
rect 511264 2926 511316 2932
rect 511276 480 511304 2926
rect 512472 480 512500 4218
rect 513576 480 513604 6122
rect 514772 480 514800 148514
rect 522304 148504 522356 148510
rect 522304 148446 522356 148452
rect 520280 147416 520332 147422
rect 520280 147358 520332 147364
rect 517152 7880 517204 7886
rect 517152 7822 517204 7828
rect 515956 4344 516008 4350
rect 515956 4286 516008 4292
rect 515968 480 515996 4286
rect 517164 480 517192 7822
rect 519544 4412 519596 4418
rect 519544 4354 519596 4360
rect 518348 3052 518400 3058
rect 518348 2994 518400 3000
rect 518360 480 518388 2994
rect 519556 480 519584 4354
rect 520292 490 520320 147358
rect 522316 4214 522344 148446
rect 526444 148436 526496 148442
rect 526444 148378 526496 148384
rect 523040 4548 523092 4554
rect 523040 4490 523092 4496
rect 522304 4208 522356 4214
rect 522304 4150 522356 4156
rect 521844 3120 521896 3126
rect 521844 3062 521896 3068
rect 520568 598 520780 626
rect 520568 490 520596 598
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 462 520596 490
rect 520752 480 520780 598
rect 521856 480 521884 3062
rect 523052 480 523080 4490
rect 526456 4214 526484 148378
rect 530584 148368 530636 148374
rect 530584 148310 530636 148316
rect 530124 4548 530176 4554
rect 530124 4490 530176 4496
rect 526628 4480 526680 4486
rect 526628 4422 526680 4428
rect 524236 4208 524288 4214
rect 524236 4150 524288 4156
rect 526444 4208 526496 4214
rect 526444 4150 526496 4156
rect 524248 480 524276 4150
rect 525432 3188 525484 3194
rect 525432 3130 525484 3136
rect 525444 480 525472 3130
rect 526640 480 526668 4422
rect 527824 4208 527876 4214
rect 527824 4150 527876 4156
rect 527836 480 527864 4150
rect 529020 3256 529072 3262
rect 529020 3198 529072 3204
rect 529032 480 529060 3198
rect 530136 480 530164 4490
rect 530596 4214 530624 148310
rect 538220 147348 538272 147354
rect 538220 147290 538272 147296
rect 538232 16574 538260 147290
rect 540244 147280 540296 147286
rect 540244 147222 540296 147228
rect 538232 16546 538444 16574
rect 534908 7812 534960 7818
rect 534908 7754 534960 7760
rect 533712 4684 533764 4690
rect 533712 4626 533764 4632
rect 530584 4208 530636 4214
rect 530584 4150 530636 4156
rect 531320 4208 531372 4214
rect 531320 4150 531372 4156
rect 531332 480 531360 4150
rect 532516 3324 532568 3330
rect 532516 3266 532568 3272
rect 532528 480 532556 3266
rect 533724 480 533752 4626
rect 534920 480 534948 7754
rect 537208 5500 537260 5506
rect 537208 5442 537260 5448
rect 536104 3392 536156 3398
rect 536104 3334 536156 3340
rect 536116 480 536144 3334
rect 537220 480 537248 5442
rect 538416 480 538444 16546
rect 539600 4140 539652 4146
rect 539600 4082 539652 4088
rect 539612 480 539640 4082
rect 540256 3398 540284 147222
rect 544384 147212 544436 147218
rect 544384 147154 544436 147160
rect 544292 5432 544344 5438
rect 544292 5374 544344 5380
rect 540796 4752 540848 4758
rect 540796 4694 540848 4700
rect 540244 3392 540296 3398
rect 540244 3334 540296 3340
rect 540808 480 540836 4694
rect 543188 4072 543240 4078
rect 543188 4014 543240 4020
rect 541992 3392 542044 3398
rect 541992 3334 542044 3340
rect 542004 480 542032 3334
rect 543200 480 543228 4014
rect 544304 2802 544332 5374
rect 544396 3398 544424 147154
rect 547880 147144 547932 147150
rect 547880 147086 547932 147092
rect 547892 16574 547920 147086
rect 551284 147076 551336 147082
rect 551284 147018 551336 147024
rect 547892 16546 548656 16574
rect 547880 5364 547932 5370
rect 547880 5306 547932 5312
rect 546684 4004 546736 4010
rect 546684 3946 546736 3952
rect 544384 3392 544436 3398
rect 544384 3334 544436 3340
rect 545488 3392 545540 3398
rect 545488 3334 545540 3340
rect 544304 2774 544424 2802
rect 544396 480 544424 2774
rect 545500 480 545528 3334
rect 546696 480 546724 3946
rect 547892 480 547920 5306
rect 548628 490 548656 16546
rect 550272 3936 550324 3942
rect 550272 3878 550324 3884
rect 548904 598 549116 626
rect 548904 490 548932 598
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 462 548932 490
rect 549088 480 549116 598
rect 550284 480 550312 3878
rect 551296 3398 551324 147018
rect 569224 147008 569276 147014
rect 569224 146950 569276 146956
rect 558184 145852 558236 145858
rect 558184 145794 558236 145800
rect 556252 145784 556304 145790
rect 556252 145726 556304 145732
rect 556264 6914 556292 145726
rect 556172 6886 556292 6914
rect 551468 5296 551520 5302
rect 551468 5238 551520 5244
rect 551284 3392 551336 3398
rect 551284 3334 551336 3340
rect 551480 480 551508 5238
rect 554964 5228 555016 5234
rect 554964 5170 555016 5176
rect 553768 3868 553820 3874
rect 553768 3810 553820 3816
rect 552664 3392 552716 3398
rect 552664 3334 552716 3340
rect 552676 480 552704 3334
rect 553780 480 553808 3810
rect 554976 480 555004 5170
rect 556172 480 556200 6886
rect 557356 3800 557408 3806
rect 557356 3742 557408 3748
rect 557368 480 557396 3742
rect 558196 3398 558224 145794
rect 560944 145716 560996 145722
rect 560944 145658 560996 145664
rect 558552 5160 558604 5166
rect 558552 5102 558604 5108
rect 558184 3392 558236 3398
rect 558184 3334 558236 3340
rect 558564 480 558592 5102
rect 560852 3732 560904 3738
rect 560852 3674 560904 3680
rect 559748 3392 559800 3398
rect 559748 3334 559800 3340
rect 559760 480 559788 3334
rect 560864 480 560892 3674
rect 560956 3398 560984 145658
rect 565820 145648 565872 145654
rect 565820 145590 565872 145596
rect 565832 16574 565860 145590
rect 565832 16546 566872 16574
rect 562048 5092 562100 5098
rect 562048 5034 562100 5040
rect 560944 3392 560996 3398
rect 560944 3334 560996 3340
rect 562060 480 562088 5034
rect 565636 5024 565688 5030
rect 565636 4966 565688 4972
rect 564440 3664 564492 3670
rect 564440 3606 564492 3612
rect 563244 3392 563296 3398
rect 563244 3334 563296 3340
rect 563256 480 563284 3334
rect 564452 480 564480 3606
rect 565648 480 565676 4966
rect 566844 480 566872 16546
rect 569132 4956 569184 4962
rect 569132 4898 569184 4904
rect 568028 3528 568080 3534
rect 568028 3470 568080 3476
rect 568040 480 568068 3470
rect 569144 480 569172 4898
rect 569236 3534 569264 146950
rect 572720 146940 572772 146946
rect 572720 146882 572772 146888
rect 572732 16574 572760 146882
rect 574744 145580 574796 145586
rect 574744 145522 574796 145528
rect 572732 16546 573496 16574
rect 572720 4820 572772 4826
rect 572720 4762 572772 4768
rect 569224 3528 569276 3534
rect 569224 3470 569276 3476
rect 570328 3528 570380 3534
rect 570328 3470 570380 3476
rect 570340 480 570368 3470
rect 571524 3460 571576 3466
rect 571524 3402 571576 3408
rect 571536 480 571564 3402
rect 572732 480 572760 4762
rect 573468 490 573496 16546
rect 574756 4146 574784 145522
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 576308 4888 576360 4894
rect 576308 4830 576360 4836
rect 574744 4140 574796 4146
rect 574744 4082 574796 4088
rect 575110 3768 575166 3777
rect 575110 3703 575166 3712
rect 573744 598 573956 626
rect 573744 490 573772 598
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573468 462 573772 490
rect 573928 480 573956 598
rect 575124 480 575152 3703
rect 576320 480 576348 4830
rect 577412 4140 577464 4146
rect 577412 4082 577464 4088
rect 577424 480 577452 4082
rect 578606 3632 578662 3641
rect 578606 3567 578662 3576
rect 582196 3596 582248 3602
rect 578620 480 578648 3567
rect 582196 3538 582248 3544
rect 580998 3496 581054 3505
rect 580998 3431 581054 3440
rect 581012 480 581040 3431
rect 582208 480 582236 3538
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3330 553832 3386 553888
rect 3238 527856 3294 527912
rect 3330 514800 3386 514856
rect 2870 462576 2926 462632
rect 3330 397432 3386 397488
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 4066 501744 4122 501800
rect 3974 475632 4030 475688
rect 3882 449520 3938 449576
rect 3790 423544 3846 423600
rect 3698 410488 3754 410544
rect 3606 371320 3662 371376
rect 3514 319232 3570 319288
rect 3514 306176 3570 306232
rect 3422 293120 3478 293176
rect 2778 267144 2834 267200
rect 3422 254088 3478 254144
rect 3422 241032 3478 241088
rect 3330 214920 3386 214976
rect 3422 201864 3478 201920
rect 3422 188808 3478 188864
rect 3238 162832 3294 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3422 111696 3478 111752
rect 3422 110608 3478 110664
rect 3422 85448 3478 85504
rect 3422 84632 3478 84688
rect 3330 59200 3386 59256
rect 3330 58520 3386 58576
rect 3330 33088 3386 33144
rect 3330 32408 3386 32464
rect 3422 20576 3478 20632
rect 3422 19352 3478 19408
rect 5262 3304 5318 3360
rect 11150 3440 11206 3496
rect 14738 3576 14794 3632
rect 20626 3712 20682 3768
rect 131670 557504 131726 557560
rect 134614 557504 134670 557560
rect 137742 557504 137798 557560
rect 140594 557504 140650 557560
rect 143354 557504 143410 557560
rect 145930 557504 145986 557560
rect 149334 557504 149390 557560
rect 152462 557504 152518 557560
rect 158350 557504 158406 557560
rect 436650 557504 436706 557560
rect 439594 557504 439650 557560
rect 443090 557504 443146 557560
rect 445758 557504 445814 557560
rect 448610 557504 448666 557560
rect 451554 557504 451610 557560
rect 454498 557504 454554 557560
rect 457442 557504 457498 557560
rect 460386 557504 460442 557560
rect 127162 3304 127218 3360
rect 129922 3440 129978 3496
rect 132590 3576 132646 3632
rect 135350 3712 135406 3768
rect 456614 3476 456616 3496
rect 456616 3476 456668 3496
rect 456668 3476 456670 3496
rect 456614 3440 456670 3476
rect 457994 3712 458050 3768
rect 458178 3476 458180 3496
rect 458180 3476 458232 3496
rect 458232 3476 458234 3496
rect 458178 3440 458234 3476
rect 460846 3576 460902 3632
rect 460754 3440 460810 3496
rect 462134 3304 462190 3360
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 580170 418240 580226 418296
rect 579618 404912 579674 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 579894 325216 579950 325272
rect 580170 312024 580226 312080
rect 579618 298696 579674 298752
rect 579894 272176 579950 272232
rect 579802 258848 579858 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 232328 580226 232384
rect 579894 219000 579950 219056
rect 580170 205672 580226 205728
rect 580170 192480 580226 192536
rect 579986 179152 580042 179208
rect 580814 537784 580870 537840
rect 580722 524456 580778 524512
rect 580630 511264 580686 511320
rect 580538 484608 580594 484664
rect 580446 471416 580502 471472
rect 580354 431568 580410 431624
rect 580262 165824 580318 165880
rect 580170 152632 580226 152688
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 6568 580226 6624
rect 575110 3712 575166 3768
rect 578606 3576 578662 3632
rect 580998 3440 581054 3496
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect 131665 557562 131731 557565
rect 132350 557562 132356 557564
rect 131665 557560 132356 557562
rect 131665 557504 131670 557560
rect 131726 557504 132356 557560
rect 131665 557502 132356 557504
rect 131665 557499 131731 557502
rect 132350 557500 132356 557502
rect 132420 557500 132426 557564
rect 134609 557562 134675 557565
rect 134926 557562 134932 557564
rect 134609 557560 134932 557562
rect 134609 557504 134614 557560
rect 134670 557504 134932 557560
rect 134609 557502 134932 557504
rect 134609 557499 134675 557502
rect 134926 557500 134932 557502
rect 134996 557500 135002 557564
rect 137737 557562 137803 557565
rect 140589 557564 140655 557565
rect 143349 557564 143415 557565
rect 137870 557562 137876 557564
rect 137737 557560 137876 557562
rect 137737 557504 137742 557560
rect 137798 557504 137876 557560
rect 137737 557502 137876 557504
rect 137737 557499 137803 557502
rect 137870 557500 137876 557502
rect 137940 557500 137946 557564
rect 140589 557560 140636 557564
rect 140700 557562 140706 557564
rect 140589 557504 140594 557560
rect 140589 557500 140636 557504
rect 140700 557502 140746 557562
rect 143349 557560 143396 557564
rect 143460 557562 143466 557564
rect 143349 557504 143354 557560
rect 140700 557500 140706 557502
rect 143349 557500 143396 557504
rect 143460 557502 143506 557562
rect 143460 557500 143466 557502
rect 145598 557500 145604 557564
rect 145668 557562 145674 557564
rect 145925 557562 145991 557565
rect 149329 557564 149395 557565
rect 149278 557562 149284 557564
rect 145668 557560 145991 557562
rect 145668 557504 145930 557560
rect 145986 557504 145991 557560
rect 145668 557502 145991 557504
rect 149238 557502 149284 557562
rect 149348 557560 149395 557564
rect 149390 557504 149395 557560
rect 145668 557500 145674 557502
rect 140589 557499 140655 557500
rect 143349 557499 143415 557500
rect 145925 557499 145991 557502
rect 149278 557500 149284 557502
rect 149348 557500 149395 557504
rect 149329 557499 149395 557500
rect 152457 557562 152523 557565
rect 152958 557562 152964 557564
rect 152457 557560 152964 557562
rect 152457 557504 152462 557560
rect 152518 557504 152964 557560
rect 152457 557502 152964 557504
rect 152457 557499 152523 557502
rect 152958 557500 152964 557502
rect 153028 557500 153034 557564
rect 158345 557562 158411 557565
rect 158478 557562 158484 557564
rect 158345 557560 158484 557562
rect 158345 557504 158350 557560
rect 158406 557504 158484 557560
rect 158345 557502 158484 557504
rect 158345 557499 158411 557502
rect 158478 557500 158484 557502
rect 158548 557500 158554 557564
rect 436134 557500 436140 557564
rect 436204 557562 436210 557564
rect 436645 557562 436711 557565
rect 436204 557560 436711 557562
rect 436204 557504 436650 557560
rect 436706 557504 436711 557560
rect 436204 557502 436711 557504
rect 436204 557500 436210 557502
rect 436645 557499 436711 557502
rect 438894 557500 438900 557564
rect 438964 557562 438970 557564
rect 439589 557562 439655 557565
rect 438964 557560 439655 557562
rect 438964 557504 439594 557560
rect 439650 557504 439655 557560
rect 438964 557502 439655 557504
rect 438964 557500 438970 557502
rect 439589 557499 439655 557502
rect 442942 557500 442948 557564
rect 443012 557562 443018 557564
rect 443085 557562 443151 557565
rect 445753 557564 445819 557565
rect 445702 557562 445708 557564
rect 443012 557560 443151 557562
rect 443012 557504 443090 557560
rect 443146 557504 443151 557560
rect 443012 557502 443151 557504
rect 445662 557502 445708 557562
rect 445772 557560 445819 557564
rect 445814 557504 445819 557560
rect 443012 557500 443018 557502
rect 443085 557499 443151 557502
rect 445702 557500 445708 557502
rect 445772 557500 445819 557504
rect 448462 557500 448468 557564
rect 448532 557562 448538 557564
rect 448605 557562 448671 557565
rect 448532 557560 448671 557562
rect 448532 557504 448610 557560
rect 448666 557504 448671 557560
rect 448532 557502 448671 557504
rect 448532 557500 448538 557502
rect 445753 557499 445819 557500
rect 448605 557499 448671 557502
rect 451222 557500 451228 557564
rect 451292 557562 451298 557564
rect 451549 557562 451615 557565
rect 451292 557560 451615 557562
rect 451292 557504 451554 557560
rect 451610 557504 451615 557560
rect 451292 557502 451615 557504
rect 451292 557500 451298 557502
rect 451549 557499 451615 557502
rect 454166 557500 454172 557564
rect 454236 557562 454242 557564
rect 454493 557562 454559 557565
rect 454236 557560 454559 557562
rect 454236 557504 454498 557560
rect 454554 557504 454559 557560
rect 454236 557502 454559 557504
rect 454236 557500 454242 557502
rect 454493 557499 454559 557502
rect 456742 557500 456748 557564
rect 456812 557562 456818 557564
rect 457437 557562 457503 557565
rect 456812 557560 457503 557562
rect 456812 557504 457442 557560
rect 457498 557504 457503 557560
rect 456812 557502 457503 557504
rect 456812 557500 456818 557502
rect 457437 557499 457503 557502
rect 460054 557500 460060 557564
rect 460124 557562 460130 557564
rect 460381 557562 460447 557565
rect 460124 557560 460447 557562
rect 460124 557504 460386 557560
rect 460442 557504 460447 557560
rect 460124 557502 460447 557504
rect 460124 557500 460130 557502
rect 460381 557499 460447 557502
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580809 537842 580875 537845
rect 583520 537842 584960 537932
rect 580809 537840 584960 537842
rect 580809 537784 580814 537840
rect 580870 537784 584960 537840
rect 580809 537782 584960 537784
rect 580809 537779 580875 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3233 527914 3299 527917
rect -960 527912 3299 527914
rect -960 527856 3238 527912
rect 3294 527856 3299 527912
rect -960 527854 3299 527856
rect -960 527764 480 527854
rect 3233 527851 3299 527854
rect 580717 524514 580783 524517
rect 583520 524514 584960 524604
rect 580717 524512 584960 524514
rect 580717 524456 580722 524512
rect 580778 524456 584960 524512
rect 580717 524454 584960 524456
rect 580717 524451 580783 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580625 511322 580691 511325
rect 583520 511322 584960 511412
rect 580625 511320 584960 511322
rect 580625 511264 580630 511320
rect 580686 511264 584960 511320
rect 580625 511262 584960 511264
rect 580625 511259 580691 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 4061 501802 4127 501805
rect -960 501800 4127 501802
rect -960 501744 4066 501800
rect 4122 501744 4127 501800
rect -960 501742 4127 501744
rect -960 501652 480 501742
rect 4061 501739 4127 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580533 484666 580599 484669
rect 583520 484666 584960 484756
rect 580533 484664 584960 484666
rect 580533 484608 580538 484664
rect 580594 484608 584960 484664
rect 580533 484606 584960 484608
rect 580533 484603 580599 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3969 475690 4035 475693
rect -960 475688 4035 475690
rect -960 475632 3974 475688
rect 4030 475632 4035 475688
rect -960 475630 4035 475632
rect -960 475540 480 475630
rect 3969 475627 4035 475630
rect 580441 471474 580507 471477
rect 583520 471474 584960 471564
rect 580441 471472 584960 471474
rect 580441 471416 580446 471472
rect 580502 471416 584960 471472
rect 580441 471414 584960 471416
rect 580441 471411 580507 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 2865 462634 2931 462637
rect -960 462632 2931 462634
rect -960 462576 2870 462632
rect 2926 462576 2931 462632
rect -960 462574 2931 462576
rect -960 462484 480 462574
rect 2865 462571 2931 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3877 449578 3943 449581
rect -960 449576 3943 449578
rect -960 449520 3882 449576
rect 3938 449520 3943 449576
rect -960 449518 3943 449520
rect -960 449428 480 449518
rect 3877 449515 3943 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580349 431626 580415 431629
rect 583520 431626 584960 431716
rect 580349 431624 584960 431626
rect 580349 431568 580354 431624
rect 580410 431568 584960 431624
rect 580349 431566 584960 431568
rect 580349 431563 580415 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3785 423602 3851 423605
rect -960 423600 3851 423602
rect -960 423544 3790 423600
rect 3846 423544 3851 423600
rect -960 423542 3851 423544
rect -960 423452 480 423542
rect 3785 423539 3851 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3693 410546 3759 410549
rect -960 410544 3759 410546
rect -960 410488 3698 410544
rect 3754 410488 3759 410544
rect -960 410486 3759 410488
rect -960 410396 480 410486
rect 3693 410483 3759 410486
rect 579613 404970 579679 404973
rect 583520 404970 584960 405060
rect 579613 404968 584960 404970
rect 579613 404912 579618 404968
rect 579674 404912 584960 404968
rect 579613 404910 584960 404912
rect 579613 404907 579679 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3601 371378 3667 371381
rect -960 371376 3667 371378
rect -960 371320 3606 371376
rect 3662 371320 3667 371376
rect -960 371318 3667 371320
rect -960 371228 480 371318
rect 3601 371315 3667 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579889 325274 579955 325277
rect 583520 325274 584960 325364
rect 579889 325272 584960 325274
rect 579889 325216 579894 325272
rect 579950 325216 584960 325272
rect 579889 325214 584960 325216
rect 579889 325211 579955 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3509 319290 3575 319293
rect -960 319288 3575 319290
rect -960 319232 3514 319288
rect 3570 319232 3575 319288
rect -960 319230 3575 319232
rect -960 319140 480 319230
rect 3509 319227 3575 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2773 267202 2839 267205
rect -960 267200 2839 267202
rect -960 267144 2778 267200
rect 2834 267144 2839 267200
rect -960 267142 2839 267144
rect -960 267052 480 267142
rect 2773 267139 2839 267142
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 579889 219058 579955 219061
rect 583520 219058 584960 219148
rect 579889 219056 584960 219058
rect 579889 219000 579894 219056
rect 579950 219000 584960 219056
rect 579889 218998 584960 219000
rect 579889 218995 579955 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 579981 179210 580047 179213
rect 583520 179210 584960 179300
rect 579981 179208 584960 179210
rect 579981 179152 579986 179208
rect 580042 179152 584960 179208
rect 579981 179150 584960 179152
rect 579981 179147 580047 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580257 165882 580323 165885
rect 583520 165882 584960 165972
rect 580257 165880 584960 165882
rect 580257 165824 580262 165880
rect 580318 165824 584960 165880
rect 580257 165822 584960 165824
rect 580257 165819 580323 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 583520 139362 584960 139452
rect 583342 139302 584960 139362
rect 583342 139226 583402 139302
rect 583520 139226 584960 139302
rect 583342 139212 584960 139226
rect 583342 139166 583586 139212
rect 158478 138076 158484 138140
rect 158548 138138 158554 138140
rect 583526 138138 583586 139166
rect 158548 138078 583586 138138
rect 158548 138076 158554 138078
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 583520 126034 584960 126124
rect 583342 125974 584960 126034
rect 583342 125898 583402 125974
rect 583520 125898 584960 125974
rect 583342 125884 584960 125898
rect 583342 125838 583586 125884
rect 152958 125564 152964 125628
rect 153028 125626 153034 125628
rect 583526 125626 583586 125838
rect 153028 125566 583586 125626
rect 153028 125564 153034 125566
rect -960 123572 480 123812
rect 583520 112842 584960 112932
rect 583342 112782 584960 112842
rect 583342 112706 583402 112782
rect 583520 112706 584960 112782
rect 583342 112692 584960 112706
rect 583342 112646 583586 112692
rect 145598 111828 145604 111892
rect 145668 111890 145674 111892
rect 583526 111890 583586 112646
rect 145668 111830 583586 111890
rect 145668 111828 145674 111830
rect 3417 111754 3483 111757
rect 436134 111754 436140 111756
rect 3417 111752 436140 111754
rect 3417 111696 3422 111752
rect 3478 111696 436140 111752
rect 3417 111694 436140 111696
rect 3417 111691 3483 111694
rect 436134 111692 436140 111694
rect 436204 111692 436210 111756
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 149278 99452 149284 99516
rect 149348 99514 149354 99516
rect 583520 99514 584960 99604
rect 149348 99454 584960 99514
rect 149348 99452 149354 99454
rect 583520 99364 584960 99454
rect 442942 97882 442948 97884
rect 6870 97822 442948 97882
rect -960 97610 480 97700
rect 6870 97610 6930 97822
rect 442942 97820 442948 97822
rect 443012 97820 443018 97884
rect -960 97550 6930 97610
rect -960 97460 480 97550
rect 583520 86186 584960 86276
rect 583342 86126 584960 86186
rect 583342 86050 583402 86126
rect 583520 86050 584960 86126
rect 583342 86036 584960 86050
rect 583342 85990 583586 86036
rect 143390 85580 143396 85644
rect 143460 85642 143466 85644
rect 583526 85642 583586 85990
rect 143460 85582 583586 85642
rect 143460 85580 143466 85582
rect 3417 85506 3483 85509
rect 438894 85506 438900 85508
rect 3417 85504 438900 85506
rect 3417 85448 3422 85504
rect 3478 85448 438900 85504
rect 3417 85446 438900 85448
rect 3417 85443 3483 85446
rect 438894 85444 438900 85446
rect 438964 85444 438970 85508
rect -960 84690 480 84780
rect 3417 84690 3483 84693
rect -960 84688 3483 84690
rect -960 84632 3422 84688
rect 3478 84632 3483 84688
rect -960 84630 3483 84632
rect -960 84540 480 84630
rect 3417 84627 3483 84630
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 137870 71844 137876 71908
rect 137940 71906 137946 71908
rect 583526 71906 583586 72798
rect 137940 71846 583586 71906
rect 137940 71844 137946 71846
rect 445702 71770 445708 71772
rect -960 71634 480 71724
rect 6870 71710 445708 71770
rect 6870 71634 6930 71710
rect 445702 71708 445708 71710
rect 445772 71708 445778 71772
rect -960 71574 6930 71634
rect -960 71484 480 71574
rect 583520 59666 584960 59756
rect 567150 59606 584960 59666
rect 140630 59332 140636 59396
rect 140700 59394 140706 59396
rect 567150 59394 567210 59606
rect 583520 59516 584960 59606
rect 140700 59334 567210 59394
rect 140700 59332 140706 59334
rect 3325 59258 3391 59261
rect 451038 59258 451044 59260
rect 3325 59256 451044 59258
rect 3325 59200 3330 59256
rect 3386 59200 451044 59256
rect 3325 59198 451044 59200
rect 3325 59195 3391 59198
rect 451038 59196 451044 59198
rect 451108 59196 451114 59260
rect -960 58578 480 58668
rect 3325 58578 3391 58581
rect -960 58576 3391 58578
rect -960 58520 3330 58576
rect 3386 58520 3391 58576
rect -960 58518 3391 58520
rect -960 58428 480 58518
rect 3325 58515 3391 58518
rect 583520 46338 584960 46428
rect 583342 46278 584960 46338
rect 583342 46202 583402 46278
rect 583520 46202 584960 46278
rect 583342 46188 584960 46202
rect 583342 46142 583586 46188
rect -960 45522 480 45612
rect 134926 45596 134932 45660
rect 134996 45658 135002 45660
rect 583526 45658 583586 46142
rect 134996 45598 583586 45658
rect 134996 45596 135002 45598
rect 448462 45522 448468 45524
rect -960 45462 448468 45522
rect -960 45372 480 45462
rect 448462 45460 448468 45462
rect 448532 45460 448538 45524
rect 3325 33146 3391 33149
rect 454166 33146 454172 33148
rect 3325 33144 454172 33146
rect 3325 33088 3330 33144
rect 3386 33088 454172 33144
rect 3325 33086 454172 33088
rect 3325 33083 3391 33086
rect 454166 33084 454172 33086
rect 454236 33084 454242 33148
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3325 32466 3391 32469
rect -960 32464 3391 32466
rect -960 32408 3330 32464
rect 3386 32408 3391 32464
rect -960 32406 3391 32408
rect -960 32316 480 32406
rect 3325 32403 3391 32406
rect 3417 20634 3483 20637
rect 460054 20634 460060 20636
rect 3417 20632 460060 20634
rect 3417 20576 3422 20632
rect 3478 20576 460060 20632
rect 3417 20574 460060 20576
rect 3417 20571 3483 20574
rect 460054 20572 460060 20574
rect 460124 20572 460130 20636
rect 583520 19818 584960 19908
rect 583342 19758 584960 19818
rect 583342 19682 583402 19758
rect 583520 19682 584960 19758
rect 583342 19668 584960 19682
rect 583342 19622 583586 19668
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 132350 19348 132356 19412
rect 132420 19410 132426 19412
rect 583526 19410 583586 19622
rect 132420 19350 583586 19410
rect 132420 19348 132426 19350
rect 456742 6898 456748 6900
rect 6870 6838 456748 6898
rect -960 6490 480 6580
rect 6870 6490 6930 6838
rect 456742 6836 456748 6838
rect 456812 6836 456818 6900
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect -960 6430 6930 6490
rect 583520 6476 584960 6566
rect -960 6340 480 6430
rect 20621 3770 20687 3773
rect 135345 3770 135411 3773
rect 20621 3768 135411 3770
rect 20621 3712 20626 3768
rect 20682 3712 135350 3768
rect 135406 3712 135411 3768
rect 20621 3710 135411 3712
rect 20621 3707 20687 3710
rect 135345 3707 135411 3710
rect 457989 3770 458055 3773
rect 575105 3770 575171 3773
rect 457989 3768 575171 3770
rect 457989 3712 457994 3768
rect 458050 3712 575110 3768
rect 575166 3712 575171 3768
rect 457989 3710 575171 3712
rect 457989 3707 458055 3710
rect 575105 3707 575171 3710
rect 14733 3634 14799 3637
rect 132585 3634 132651 3637
rect 14733 3632 132651 3634
rect 14733 3576 14738 3632
rect 14794 3576 132590 3632
rect 132646 3576 132651 3632
rect 14733 3574 132651 3576
rect 14733 3571 14799 3574
rect 132585 3571 132651 3574
rect 460841 3634 460907 3637
rect 578601 3634 578667 3637
rect 460841 3632 578667 3634
rect 460841 3576 460846 3632
rect 460902 3576 578606 3632
rect 578662 3576 578667 3632
rect 460841 3574 578667 3576
rect 460841 3571 460907 3574
rect 578601 3571 578667 3574
rect 11145 3498 11211 3501
rect 129917 3498 129983 3501
rect 11145 3496 129983 3498
rect 11145 3440 11150 3496
rect 11206 3440 129922 3496
rect 129978 3440 129983 3496
rect 11145 3438 129983 3440
rect 11145 3435 11211 3438
rect 129917 3435 129983 3438
rect 456609 3498 456675 3501
rect 458173 3498 458239 3501
rect 456609 3496 458239 3498
rect 456609 3440 456614 3496
rect 456670 3440 458178 3496
rect 458234 3440 458239 3496
rect 456609 3438 458239 3440
rect 456609 3435 456675 3438
rect 458173 3435 458239 3438
rect 460749 3498 460815 3501
rect 580993 3498 581059 3501
rect 460749 3496 581059 3498
rect 460749 3440 460754 3496
rect 460810 3440 580998 3496
rect 581054 3440 581059 3496
rect 460749 3438 581059 3440
rect 460749 3435 460815 3438
rect 580993 3435 581059 3438
rect 5257 3362 5323 3365
rect 127157 3362 127223 3365
rect 5257 3360 127223 3362
rect 5257 3304 5262 3360
rect 5318 3304 127162 3360
rect 127218 3304 127223 3360
rect 5257 3302 127223 3304
rect 5257 3299 5323 3302
rect 127157 3299 127223 3302
rect 462129 3362 462195 3365
rect 583385 3362 583451 3365
rect 462129 3360 583451 3362
rect 462129 3304 462134 3360
rect 462190 3304 583390 3360
rect 583446 3304 583451 3360
rect 462129 3302 583451 3304
rect 462129 3299 462195 3302
rect 583385 3299 583451 3302
<< via3 >>
rect 132356 557500 132420 557564
rect 134932 557500 134996 557564
rect 137876 557500 137940 557564
rect 140636 557560 140700 557564
rect 140636 557504 140650 557560
rect 140650 557504 140700 557560
rect 140636 557500 140700 557504
rect 143396 557560 143460 557564
rect 143396 557504 143410 557560
rect 143410 557504 143460 557560
rect 143396 557500 143460 557504
rect 145604 557500 145668 557564
rect 149284 557560 149348 557564
rect 149284 557504 149334 557560
rect 149334 557504 149348 557560
rect 149284 557500 149348 557504
rect 152964 557500 153028 557564
rect 158484 557500 158548 557564
rect 436140 557500 436204 557564
rect 438900 557500 438964 557564
rect 442948 557500 443012 557564
rect 445708 557560 445772 557564
rect 445708 557504 445758 557560
rect 445758 557504 445772 557560
rect 445708 557500 445772 557504
rect 448468 557500 448532 557564
rect 451228 557500 451292 557564
rect 454172 557500 454236 557564
rect 456748 557500 456812 557564
rect 460060 557500 460124 557564
rect 158484 138076 158548 138140
rect 152964 125564 153028 125628
rect 145604 111828 145668 111892
rect 436140 111692 436204 111756
rect 149284 99452 149348 99516
rect 442948 97820 443012 97884
rect 143396 85580 143460 85644
rect 438900 85444 438964 85508
rect 137876 71844 137940 71908
rect 445708 71708 445772 71772
rect 140636 59332 140700 59396
rect 451044 59196 451108 59260
rect 134932 45596 134996 45660
rect 448468 45460 448532 45524
rect 454172 33084 454236 33148
rect 460060 20572 460124 20636
rect 132356 19348 132420 19412
rect 456748 6836 456812 6900
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 560023 128414 560898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 560023 132134 564618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 560023 135854 568338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 560023 139574 572058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 560023 146414 578898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 560023 150134 582618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 560023 153854 586338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 560023 157574 590058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 560023 164414 560898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 560023 168134 564618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 560023 171854 568338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 560023 175574 572058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 560023 182414 578898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 560023 186134 582618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 560023 189854 586338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 560023 193574 590058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 560023 200414 560898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 560023 204134 564618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 560023 207854 568338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 560023 211574 572058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 560023 218414 578898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 560023 222134 582618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 560023 225854 586338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 560023 229574 590058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 560023 236414 560898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 560023 240134 564618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 560023 243854 568338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 560023 247574 572058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 560023 254414 578898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 560023 258134 582618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 560023 261854 586338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 560023 265574 590058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 560023 272414 560898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 560023 276134 564618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 560023 279854 568338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 560023 283574 572058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 560023 290414 578898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 560023 294134 582618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 560023 297854 586338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 560023 301574 590058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 560023 308414 560898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 560023 312134 564618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 560023 315854 568338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 560023 319574 572058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 560023 326414 578898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 560023 330134 582618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 560023 333854 586338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 560023 337574 590058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 560023 344414 560898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 560023 348134 564618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 560023 351854 568338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 560023 355574 572058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 560023 362414 578898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 560023 366134 582618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 560023 369854 586338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 560023 373574 590058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 560023 380414 560898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 560023 384134 564618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 560023 387854 568338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 560023 391574 572058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 560023 398414 578898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 560023 402134 582618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 560023 405854 586338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 560023 409574 590058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 560023 416414 560898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 560023 420134 564618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 560023 423854 568338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 560023 427574 572058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 560023 434414 578898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 560023 438134 582618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 560023 441854 586338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 560023 445574 590058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 560023 452414 560898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 560023 456134 564618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 560023 459854 568338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 560023 463574 572058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 132355 557564 132421 557565
rect 132355 557500 132356 557564
rect 132420 557500 132421 557564
rect 132355 557499 132421 557500
rect 134931 557564 134997 557565
rect 134931 557500 134932 557564
rect 134996 557500 134997 557564
rect 134931 557499 134997 557500
rect 137875 557564 137941 557565
rect 137875 557500 137876 557564
rect 137940 557500 137941 557564
rect 137875 557499 137941 557500
rect 140635 557564 140701 557565
rect 140635 557500 140636 557564
rect 140700 557500 140701 557564
rect 140635 557499 140701 557500
rect 143395 557564 143461 557565
rect 143395 557500 143396 557564
rect 143460 557500 143461 557564
rect 143395 557499 143461 557500
rect 145603 557564 145669 557565
rect 145603 557500 145604 557564
rect 145668 557500 145669 557564
rect 145603 557499 145669 557500
rect 149283 557564 149349 557565
rect 149283 557500 149284 557564
rect 149348 557500 149349 557564
rect 149283 557499 149349 557500
rect 152963 557564 153029 557565
rect 152963 557500 152964 557564
rect 153028 557500 153029 557564
rect 152963 557499 153029 557500
rect 158483 557564 158549 557565
rect 158483 557500 158484 557564
rect 158548 557500 158549 557564
rect 158483 557499 158549 557500
rect 436139 557564 436205 557565
rect 436139 557500 436140 557564
rect 436204 557500 436205 557564
rect 436139 557499 436205 557500
rect 438899 557564 438965 557565
rect 438899 557500 438900 557564
rect 438964 557500 438965 557564
rect 438899 557499 438965 557500
rect 442947 557564 443013 557565
rect 442947 557500 442948 557564
rect 443012 557500 443013 557564
rect 442947 557499 443013 557500
rect 445707 557564 445773 557565
rect 445707 557500 445708 557564
rect 445772 557500 445773 557564
rect 445707 557499 445773 557500
rect 448467 557564 448533 557565
rect 448467 557500 448468 557564
rect 448532 557500 448533 557564
rect 451227 557564 451293 557565
rect 451227 557550 451228 557564
rect 448467 557499 448533 557500
rect 451046 557500 451228 557550
rect 451292 557500 451293 557564
rect 451046 557499 451293 557500
rect 454171 557564 454237 557565
rect 454171 557500 454172 557564
rect 454236 557500 454237 557564
rect 454171 557499 454237 557500
rect 456747 557564 456813 557565
rect 456747 557500 456748 557564
rect 456812 557500 456813 557564
rect 456747 557499 456813 557500
rect 460059 557564 460125 557565
rect 460059 557500 460060 557564
rect 460124 557500 460125 557564
rect 460059 557499 460125 557500
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 128208 543454 128528 543486
rect 128208 543218 128250 543454
rect 128486 543218 128528 543454
rect 128208 543134 128528 543218
rect 128208 542898 128250 543134
rect 128486 542898 128528 543134
rect 128208 542866 128528 542898
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 128208 507454 128528 507486
rect 128208 507218 128250 507454
rect 128486 507218 128528 507454
rect 128208 507134 128528 507218
rect 128208 506898 128250 507134
rect 128486 506898 128528 507134
rect 128208 506866 128528 506898
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 128208 471454 128528 471486
rect 128208 471218 128250 471454
rect 128486 471218 128528 471454
rect 128208 471134 128528 471218
rect 128208 470898 128250 471134
rect 128486 470898 128528 471134
rect 128208 470866 128528 470898
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 128208 435454 128528 435486
rect 128208 435218 128250 435454
rect 128486 435218 128528 435454
rect 128208 435134 128528 435218
rect 128208 434898 128250 435134
rect 128486 434898 128528 435134
rect 128208 434866 128528 434898
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 128208 399454 128528 399486
rect 128208 399218 128250 399454
rect 128486 399218 128528 399454
rect 128208 399134 128528 399218
rect 128208 398898 128250 399134
rect 128486 398898 128528 399134
rect 128208 398866 128528 398898
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 128208 363454 128528 363486
rect 128208 363218 128250 363454
rect 128486 363218 128528 363454
rect 128208 363134 128528 363218
rect 128208 362898 128250 363134
rect 128486 362898 128528 363134
rect 128208 362866 128528 362898
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 128208 327454 128528 327486
rect 128208 327218 128250 327454
rect 128486 327218 128528 327454
rect 128208 327134 128528 327218
rect 128208 326898 128250 327134
rect 128486 326898 128528 327134
rect 128208 326866 128528 326898
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 128208 291454 128528 291486
rect 128208 291218 128250 291454
rect 128486 291218 128528 291454
rect 128208 291134 128528 291218
rect 128208 290898 128250 291134
rect 128486 290898 128528 291134
rect 128208 290866 128528 290898
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 128208 255454 128528 255486
rect 128208 255218 128250 255454
rect 128486 255218 128528 255454
rect 128208 255134 128528 255218
rect 128208 254898 128250 255134
rect 128486 254898 128528 255134
rect 128208 254866 128528 254898
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 128208 219454 128528 219486
rect 128208 219218 128250 219454
rect 128486 219218 128528 219454
rect 128208 219134 128528 219218
rect 128208 218898 128250 219134
rect 128486 218898 128528 219134
rect 128208 218866 128528 218898
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 128208 183454 128528 183486
rect 128208 183218 128250 183454
rect 128486 183218 128528 183454
rect 128208 183134 128528 183218
rect 128208 182898 128250 183134
rect 128486 182898 128528 183134
rect 128208 182866 128528 182898
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 129454 128414 148400
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 133174 132134 148400
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 132358 19413 132418 557499
rect 134934 45661 134994 557499
rect 135234 136894 135854 148400
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 137878 71909 137938 557499
rect 138954 140614 139574 148400
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 137875 71908 137941 71909
rect 137875 71844 137876 71908
rect 137940 71844 137941 71908
rect 137875 71843 137941 71844
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 134931 45660 134997 45661
rect 134931 45596 134932 45660
rect 134996 45596 134997 45660
rect 134931 45595 134997 45596
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 132355 19412 132421 19413
rect 132355 19348 132356 19412
rect 132420 19348 132421 19412
rect 132355 19347 132421 19348
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 140638 59397 140698 557499
rect 143398 85645 143458 557499
rect 143568 525454 143888 525486
rect 143568 525218 143610 525454
rect 143846 525218 143888 525454
rect 143568 525134 143888 525218
rect 143568 524898 143610 525134
rect 143846 524898 143888 525134
rect 143568 524866 143888 524898
rect 143568 489454 143888 489486
rect 143568 489218 143610 489454
rect 143846 489218 143888 489454
rect 143568 489134 143888 489218
rect 143568 488898 143610 489134
rect 143846 488898 143888 489134
rect 143568 488866 143888 488898
rect 143568 453454 143888 453486
rect 143568 453218 143610 453454
rect 143846 453218 143888 453454
rect 143568 453134 143888 453218
rect 143568 452898 143610 453134
rect 143846 452898 143888 453134
rect 143568 452866 143888 452898
rect 143568 417454 143888 417486
rect 143568 417218 143610 417454
rect 143846 417218 143888 417454
rect 143568 417134 143888 417218
rect 143568 416898 143610 417134
rect 143846 416898 143888 417134
rect 143568 416866 143888 416898
rect 143568 381454 143888 381486
rect 143568 381218 143610 381454
rect 143846 381218 143888 381454
rect 143568 381134 143888 381218
rect 143568 380898 143610 381134
rect 143846 380898 143888 381134
rect 143568 380866 143888 380898
rect 143568 345454 143888 345486
rect 143568 345218 143610 345454
rect 143846 345218 143888 345454
rect 143568 345134 143888 345218
rect 143568 344898 143610 345134
rect 143846 344898 143888 345134
rect 143568 344866 143888 344898
rect 143568 309454 143888 309486
rect 143568 309218 143610 309454
rect 143846 309218 143888 309454
rect 143568 309134 143888 309218
rect 143568 308898 143610 309134
rect 143846 308898 143888 309134
rect 143568 308866 143888 308898
rect 143568 273454 143888 273486
rect 143568 273218 143610 273454
rect 143846 273218 143888 273454
rect 143568 273134 143888 273218
rect 143568 272898 143610 273134
rect 143846 272898 143888 273134
rect 143568 272866 143888 272898
rect 143568 237454 143888 237486
rect 143568 237218 143610 237454
rect 143846 237218 143888 237454
rect 143568 237134 143888 237218
rect 143568 236898 143610 237134
rect 143846 236898 143888 237134
rect 143568 236866 143888 236898
rect 143568 201454 143888 201486
rect 143568 201218 143610 201454
rect 143846 201218 143888 201454
rect 143568 201134 143888 201218
rect 143568 200898 143610 201134
rect 143846 200898 143888 201134
rect 143568 200866 143888 200898
rect 143568 165454 143888 165486
rect 143568 165218 143610 165454
rect 143846 165218 143888 165454
rect 143568 165134 143888 165218
rect 143568 164898 143610 165134
rect 143846 164898 143888 165134
rect 143568 164866 143888 164898
rect 145606 111893 145666 557499
rect 145794 147454 146414 148400
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145603 111892 145669 111893
rect 145603 111828 145604 111892
rect 145668 111828 145669 111892
rect 145603 111827 145669 111828
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 143395 85644 143461 85645
rect 143395 85580 143396 85644
rect 143460 85580 143461 85644
rect 143395 85579 143461 85580
rect 145794 75454 146414 110898
rect 149286 99517 149346 557499
rect 149514 115174 150134 148400
rect 152966 125629 153026 557499
rect 152963 125628 153029 125629
rect 152963 125564 152964 125628
rect 153028 125564 153029 125628
rect 152963 125563 153029 125564
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149283 99516 149349 99517
rect 149283 99452 149284 99516
rect 149348 99452 149349 99516
rect 149283 99451 149349 99452
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 140635 59396 140701 59397
rect 140635 59332 140636 59396
rect 140700 59332 140701 59396
rect 140635 59331 140701 59332
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 118894 153854 148400
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 122614 157574 148400
rect 158486 138141 158546 557499
rect 158928 543454 159248 543486
rect 158928 543218 158970 543454
rect 159206 543218 159248 543454
rect 158928 543134 159248 543218
rect 158928 542898 158970 543134
rect 159206 542898 159248 543134
rect 158928 542866 159248 542898
rect 189648 543454 189968 543486
rect 189648 543218 189690 543454
rect 189926 543218 189968 543454
rect 189648 543134 189968 543218
rect 189648 542898 189690 543134
rect 189926 542898 189968 543134
rect 189648 542866 189968 542898
rect 220368 543454 220688 543486
rect 220368 543218 220410 543454
rect 220646 543218 220688 543454
rect 220368 543134 220688 543218
rect 220368 542898 220410 543134
rect 220646 542898 220688 543134
rect 220368 542866 220688 542898
rect 251088 543454 251408 543486
rect 251088 543218 251130 543454
rect 251366 543218 251408 543454
rect 251088 543134 251408 543218
rect 251088 542898 251130 543134
rect 251366 542898 251408 543134
rect 251088 542866 251408 542898
rect 281808 543454 282128 543486
rect 281808 543218 281850 543454
rect 282086 543218 282128 543454
rect 281808 543134 282128 543218
rect 281808 542898 281850 543134
rect 282086 542898 282128 543134
rect 281808 542866 282128 542898
rect 312528 543454 312848 543486
rect 312528 543218 312570 543454
rect 312806 543218 312848 543454
rect 312528 543134 312848 543218
rect 312528 542898 312570 543134
rect 312806 542898 312848 543134
rect 312528 542866 312848 542898
rect 343248 543454 343568 543486
rect 343248 543218 343290 543454
rect 343526 543218 343568 543454
rect 343248 543134 343568 543218
rect 343248 542898 343290 543134
rect 343526 542898 343568 543134
rect 343248 542866 343568 542898
rect 373968 543454 374288 543486
rect 373968 543218 374010 543454
rect 374246 543218 374288 543454
rect 373968 543134 374288 543218
rect 373968 542898 374010 543134
rect 374246 542898 374288 543134
rect 373968 542866 374288 542898
rect 404688 543454 405008 543486
rect 404688 543218 404730 543454
rect 404966 543218 405008 543454
rect 404688 543134 405008 543218
rect 404688 542898 404730 543134
rect 404966 542898 405008 543134
rect 404688 542866 405008 542898
rect 435408 543454 435728 543486
rect 435408 543218 435450 543454
rect 435686 543218 435728 543454
rect 435408 543134 435728 543218
rect 435408 542898 435450 543134
rect 435686 542898 435728 543134
rect 435408 542866 435728 542898
rect 174288 525454 174608 525486
rect 174288 525218 174330 525454
rect 174566 525218 174608 525454
rect 174288 525134 174608 525218
rect 174288 524898 174330 525134
rect 174566 524898 174608 525134
rect 174288 524866 174608 524898
rect 205008 525454 205328 525486
rect 205008 525218 205050 525454
rect 205286 525218 205328 525454
rect 205008 525134 205328 525218
rect 205008 524898 205050 525134
rect 205286 524898 205328 525134
rect 205008 524866 205328 524898
rect 235728 525454 236048 525486
rect 235728 525218 235770 525454
rect 236006 525218 236048 525454
rect 235728 525134 236048 525218
rect 235728 524898 235770 525134
rect 236006 524898 236048 525134
rect 235728 524866 236048 524898
rect 266448 525454 266768 525486
rect 266448 525218 266490 525454
rect 266726 525218 266768 525454
rect 266448 525134 266768 525218
rect 266448 524898 266490 525134
rect 266726 524898 266768 525134
rect 266448 524866 266768 524898
rect 297168 525454 297488 525486
rect 297168 525218 297210 525454
rect 297446 525218 297488 525454
rect 297168 525134 297488 525218
rect 297168 524898 297210 525134
rect 297446 524898 297488 525134
rect 297168 524866 297488 524898
rect 327888 525454 328208 525486
rect 327888 525218 327930 525454
rect 328166 525218 328208 525454
rect 327888 525134 328208 525218
rect 327888 524898 327930 525134
rect 328166 524898 328208 525134
rect 327888 524866 328208 524898
rect 358608 525454 358928 525486
rect 358608 525218 358650 525454
rect 358886 525218 358928 525454
rect 358608 525134 358928 525218
rect 358608 524898 358650 525134
rect 358886 524898 358928 525134
rect 358608 524866 358928 524898
rect 389328 525454 389648 525486
rect 389328 525218 389370 525454
rect 389606 525218 389648 525454
rect 389328 525134 389648 525218
rect 389328 524898 389370 525134
rect 389606 524898 389648 525134
rect 389328 524866 389648 524898
rect 420048 525454 420368 525486
rect 420048 525218 420090 525454
rect 420326 525218 420368 525454
rect 420048 525134 420368 525218
rect 420048 524898 420090 525134
rect 420326 524898 420368 525134
rect 420048 524866 420368 524898
rect 158928 507454 159248 507486
rect 158928 507218 158970 507454
rect 159206 507218 159248 507454
rect 158928 507134 159248 507218
rect 158928 506898 158970 507134
rect 159206 506898 159248 507134
rect 158928 506866 159248 506898
rect 189648 507454 189968 507486
rect 189648 507218 189690 507454
rect 189926 507218 189968 507454
rect 189648 507134 189968 507218
rect 189648 506898 189690 507134
rect 189926 506898 189968 507134
rect 189648 506866 189968 506898
rect 220368 507454 220688 507486
rect 220368 507218 220410 507454
rect 220646 507218 220688 507454
rect 220368 507134 220688 507218
rect 220368 506898 220410 507134
rect 220646 506898 220688 507134
rect 220368 506866 220688 506898
rect 251088 507454 251408 507486
rect 251088 507218 251130 507454
rect 251366 507218 251408 507454
rect 251088 507134 251408 507218
rect 251088 506898 251130 507134
rect 251366 506898 251408 507134
rect 251088 506866 251408 506898
rect 281808 507454 282128 507486
rect 281808 507218 281850 507454
rect 282086 507218 282128 507454
rect 281808 507134 282128 507218
rect 281808 506898 281850 507134
rect 282086 506898 282128 507134
rect 281808 506866 282128 506898
rect 312528 507454 312848 507486
rect 312528 507218 312570 507454
rect 312806 507218 312848 507454
rect 312528 507134 312848 507218
rect 312528 506898 312570 507134
rect 312806 506898 312848 507134
rect 312528 506866 312848 506898
rect 343248 507454 343568 507486
rect 343248 507218 343290 507454
rect 343526 507218 343568 507454
rect 343248 507134 343568 507218
rect 343248 506898 343290 507134
rect 343526 506898 343568 507134
rect 343248 506866 343568 506898
rect 373968 507454 374288 507486
rect 373968 507218 374010 507454
rect 374246 507218 374288 507454
rect 373968 507134 374288 507218
rect 373968 506898 374010 507134
rect 374246 506898 374288 507134
rect 373968 506866 374288 506898
rect 404688 507454 405008 507486
rect 404688 507218 404730 507454
rect 404966 507218 405008 507454
rect 404688 507134 405008 507218
rect 404688 506898 404730 507134
rect 404966 506898 405008 507134
rect 404688 506866 405008 506898
rect 435408 507454 435728 507486
rect 435408 507218 435450 507454
rect 435686 507218 435728 507454
rect 435408 507134 435728 507218
rect 435408 506898 435450 507134
rect 435686 506898 435728 507134
rect 435408 506866 435728 506898
rect 174288 489454 174608 489486
rect 174288 489218 174330 489454
rect 174566 489218 174608 489454
rect 174288 489134 174608 489218
rect 174288 488898 174330 489134
rect 174566 488898 174608 489134
rect 174288 488866 174608 488898
rect 205008 489454 205328 489486
rect 205008 489218 205050 489454
rect 205286 489218 205328 489454
rect 205008 489134 205328 489218
rect 205008 488898 205050 489134
rect 205286 488898 205328 489134
rect 205008 488866 205328 488898
rect 235728 489454 236048 489486
rect 235728 489218 235770 489454
rect 236006 489218 236048 489454
rect 235728 489134 236048 489218
rect 235728 488898 235770 489134
rect 236006 488898 236048 489134
rect 235728 488866 236048 488898
rect 266448 489454 266768 489486
rect 266448 489218 266490 489454
rect 266726 489218 266768 489454
rect 266448 489134 266768 489218
rect 266448 488898 266490 489134
rect 266726 488898 266768 489134
rect 266448 488866 266768 488898
rect 297168 489454 297488 489486
rect 297168 489218 297210 489454
rect 297446 489218 297488 489454
rect 297168 489134 297488 489218
rect 297168 488898 297210 489134
rect 297446 488898 297488 489134
rect 297168 488866 297488 488898
rect 327888 489454 328208 489486
rect 327888 489218 327930 489454
rect 328166 489218 328208 489454
rect 327888 489134 328208 489218
rect 327888 488898 327930 489134
rect 328166 488898 328208 489134
rect 327888 488866 328208 488898
rect 358608 489454 358928 489486
rect 358608 489218 358650 489454
rect 358886 489218 358928 489454
rect 358608 489134 358928 489218
rect 358608 488898 358650 489134
rect 358886 488898 358928 489134
rect 358608 488866 358928 488898
rect 389328 489454 389648 489486
rect 389328 489218 389370 489454
rect 389606 489218 389648 489454
rect 389328 489134 389648 489218
rect 389328 488898 389370 489134
rect 389606 488898 389648 489134
rect 389328 488866 389648 488898
rect 420048 489454 420368 489486
rect 420048 489218 420090 489454
rect 420326 489218 420368 489454
rect 420048 489134 420368 489218
rect 420048 488898 420090 489134
rect 420326 488898 420368 489134
rect 420048 488866 420368 488898
rect 158928 471454 159248 471486
rect 158928 471218 158970 471454
rect 159206 471218 159248 471454
rect 158928 471134 159248 471218
rect 158928 470898 158970 471134
rect 159206 470898 159248 471134
rect 158928 470866 159248 470898
rect 189648 471454 189968 471486
rect 189648 471218 189690 471454
rect 189926 471218 189968 471454
rect 189648 471134 189968 471218
rect 189648 470898 189690 471134
rect 189926 470898 189968 471134
rect 189648 470866 189968 470898
rect 220368 471454 220688 471486
rect 220368 471218 220410 471454
rect 220646 471218 220688 471454
rect 220368 471134 220688 471218
rect 220368 470898 220410 471134
rect 220646 470898 220688 471134
rect 220368 470866 220688 470898
rect 251088 471454 251408 471486
rect 251088 471218 251130 471454
rect 251366 471218 251408 471454
rect 251088 471134 251408 471218
rect 251088 470898 251130 471134
rect 251366 470898 251408 471134
rect 251088 470866 251408 470898
rect 281808 471454 282128 471486
rect 281808 471218 281850 471454
rect 282086 471218 282128 471454
rect 281808 471134 282128 471218
rect 281808 470898 281850 471134
rect 282086 470898 282128 471134
rect 281808 470866 282128 470898
rect 312528 471454 312848 471486
rect 312528 471218 312570 471454
rect 312806 471218 312848 471454
rect 312528 471134 312848 471218
rect 312528 470898 312570 471134
rect 312806 470898 312848 471134
rect 312528 470866 312848 470898
rect 343248 471454 343568 471486
rect 343248 471218 343290 471454
rect 343526 471218 343568 471454
rect 343248 471134 343568 471218
rect 343248 470898 343290 471134
rect 343526 470898 343568 471134
rect 343248 470866 343568 470898
rect 373968 471454 374288 471486
rect 373968 471218 374010 471454
rect 374246 471218 374288 471454
rect 373968 471134 374288 471218
rect 373968 470898 374010 471134
rect 374246 470898 374288 471134
rect 373968 470866 374288 470898
rect 404688 471454 405008 471486
rect 404688 471218 404730 471454
rect 404966 471218 405008 471454
rect 404688 471134 405008 471218
rect 404688 470898 404730 471134
rect 404966 470898 405008 471134
rect 404688 470866 405008 470898
rect 435408 471454 435728 471486
rect 435408 471218 435450 471454
rect 435686 471218 435728 471454
rect 435408 471134 435728 471218
rect 435408 470898 435450 471134
rect 435686 470898 435728 471134
rect 435408 470866 435728 470898
rect 174288 453454 174608 453486
rect 174288 453218 174330 453454
rect 174566 453218 174608 453454
rect 174288 453134 174608 453218
rect 174288 452898 174330 453134
rect 174566 452898 174608 453134
rect 174288 452866 174608 452898
rect 205008 453454 205328 453486
rect 205008 453218 205050 453454
rect 205286 453218 205328 453454
rect 205008 453134 205328 453218
rect 205008 452898 205050 453134
rect 205286 452898 205328 453134
rect 205008 452866 205328 452898
rect 235728 453454 236048 453486
rect 235728 453218 235770 453454
rect 236006 453218 236048 453454
rect 235728 453134 236048 453218
rect 235728 452898 235770 453134
rect 236006 452898 236048 453134
rect 235728 452866 236048 452898
rect 266448 453454 266768 453486
rect 266448 453218 266490 453454
rect 266726 453218 266768 453454
rect 266448 453134 266768 453218
rect 266448 452898 266490 453134
rect 266726 452898 266768 453134
rect 266448 452866 266768 452898
rect 297168 453454 297488 453486
rect 297168 453218 297210 453454
rect 297446 453218 297488 453454
rect 297168 453134 297488 453218
rect 297168 452898 297210 453134
rect 297446 452898 297488 453134
rect 297168 452866 297488 452898
rect 327888 453454 328208 453486
rect 327888 453218 327930 453454
rect 328166 453218 328208 453454
rect 327888 453134 328208 453218
rect 327888 452898 327930 453134
rect 328166 452898 328208 453134
rect 327888 452866 328208 452898
rect 358608 453454 358928 453486
rect 358608 453218 358650 453454
rect 358886 453218 358928 453454
rect 358608 453134 358928 453218
rect 358608 452898 358650 453134
rect 358886 452898 358928 453134
rect 358608 452866 358928 452898
rect 389328 453454 389648 453486
rect 389328 453218 389370 453454
rect 389606 453218 389648 453454
rect 389328 453134 389648 453218
rect 389328 452898 389370 453134
rect 389606 452898 389648 453134
rect 389328 452866 389648 452898
rect 420048 453454 420368 453486
rect 420048 453218 420090 453454
rect 420326 453218 420368 453454
rect 420048 453134 420368 453218
rect 420048 452898 420090 453134
rect 420326 452898 420368 453134
rect 420048 452866 420368 452898
rect 158928 435454 159248 435486
rect 158928 435218 158970 435454
rect 159206 435218 159248 435454
rect 158928 435134 159248 435218
rect 158928 434898 158970 435134
rect 159206 434898 159248 435134
rect 158928 434866 159248 434898
rect 189648 435454 189968 435486
rect 189648 435218 189690 435454
rect 189926 435218 189968 435454
rect 189648 435134 189968 435218
rect 189648 434898 189690 435134
rect 189926 434898 189968 435134
rect 189648 434866 189968 434898
rect 220368 435454 220688 435486
rect 220368 435218 220410 435454
rect 220646 435218 220688 435454
rect 220368 435134 220688 435218
rect 220368 434898 220410 435134
rect 220646 434898 220688 435134
rect 220368 434866 220688 434898
rect 251088 435454 251408 435486
rect 251088 435218 251130 435454
rect 251366 435218 251408 435454
rect 251088 435134 251408 435218
rect 251088 434898 251130 435134
rect 251366 434898 251408 435134
rect 251088 434866 251408 434898
rect 281808 435454 282128 435486
rect 281808 435218 281850 435454
rect 282086 435218 282128 435454
rect 281808 435134 282128 435218
rect 281808 434898 281850 435134
rect 282086 434898 282128 435134
rect 281808 434866 282128 434898
rect 312528 435454 312848 435486
rect 312528 435218 312570 435454
rect 312806 435218 312848 435454
rect 312528 435134 312848 435218
rect 312528 434898 312570 435134
rect 312806 434898 312848 435134
rect 312528 434866 312848 434898
rect 343248 435454 343568 435486
rect 343248 435218 343290 435454
rect 343526 435218 343568 435454
rect 343248 435134 343568 435218
rect 343248 434898 343290 435134
rect 343526 434898 343568 435134
rect 343248 434866 343568 434898
rect 373968 435454 374288 435486
rect 373968 435218 374010 435454
rect 374246 435218 374288 435454
rect 373968 435134 374288 435218
rect 373968 434898 374010 435134
rect 374246 434898 374288 435134
rect 373968 434866 374288 434898
rect 404688 435454 405008 435486
rect 404688 435218 404730 435454
rect 404966 435218 405008 435454
rect 404688 435134 405008 435218
rect 404688 434898 404730 435134
rect 404966 434898 405008 435134
rect 404688 434866 405008 434898
rect 435408 435454 435728 435486
rect 435408 435218 435450 435454
rect 435686 435218 435728 435454
rect 435408 435134 435728 435218
rect 435408 434898 435450 435134
rect 435686 434898 435728 435134
rect 435408 434866 435728 434898
rect 174288 417454 174608 417486
rect 174288 417218 174330 417454
rect 174566 417218 174608 417454
rect 174288 417134 174608 417218
rect 174288 416898 174330 417134
rect 174566 416898 174608 417134
rect 174288 416866 174608 416898
rect 205008 417454 205328 417486
rect 205008 417218 205050 417454
rect 205286 417218 205328 417454
rect 205008 417134 205328 417218
rect 205008 416898 205050 417134
rect 205286 416898 205328 417134
rect 205008 416866 205328 416898
rect 235728 417454 236048 417486
rect 235728 417218 235770 417454
rect 236006 417218 236048 417454
rect 235728 417134 236048 417218
rect 235728 416898 235770 417134
rect 236006 416898 236048 417134
rect 235728 416866 236048 416898
rect 266448 417454 266768 417486
rect 266448 417218 266490 417454
rect 266726 417218 266768 417454
rect 266448 417134 266768 417218
rect 266448 416898 266490 417134
rect 266726 416898 266768 417134
rect 266448 416866 266768 416898
rect 297168 417454 297488 417486
rect 297168 417218 297210 417454
rect 297446 417218 297488 417454
rect 297168 417134 297488 417218
rect 297168 416898 297210 417134
rect 297446 416898 297488 417134
rect 297168 416866 297488 416898
rect 327888 417454 328208 417486
rect 327888 417218 327930 417454
rect 328166 417218 328208 417454
rect 327888 417134 328208 417218
rect 327888 416898 327930 417134
rect 328166 416898 328208 417134
rect 327888 416866 328208 416898
rect 358608 417454 358928 417486
rect 358608 417218 358650 417454
rect 358886 417218 358928 417454
rect 358608 417134 358928 417218
rect 358608 416898 358650 417134
rect 358886 416898 358928 417134
rect 358608 416866 358928 416898
rect 389328 417454 389648 417486
rect 389328 417218 389370 417454
rect 389606 417218 389648 417454
rect 389328 417134 389648 417218
rect 389328 416898 389370 417134
rect 389606 416898 389648 417134
rect 389328 416866 389648 416898
rect 420048 417454 420368 417486
rect 420048 417218 420090 417454
rect 420326 417218 420368 417454
rect 420048 417134 420368 417218
rect 420048 416898 420090 417134
rect 420326 416898 420368 417134
rect 420048 416866 420368 416898
rect 158928 399454 159248 399486
rect 158928 399218 158970 399454
rect 159206 399218 159248 399454
rect 158928 399134 159248 399218
rect 158928 398898 158970 399134
rect 159206 398898 159248 399134
rect 158928 398866 159248 398898
rect 189648 399454 189968 399486
rect 189648 399218 189690 399454
rect 189926 399218 189968 399454
rect 189648 399134 189968 399218
rect 189648 398898 189690 399134
rect 189926 398898 189968 399134
rect 189648 398866 189968 398898
rect 220368 399454 220688 399486
rect 220368 399218 220410 399454
rect 220646 399218 220688 399454
rect 220368 399134 220688 399218
rect 220368 398898 220410 399134
rect 220646 398898 220688 399134
rect 220368 398866 220688 398898
rect 251088 399454 251408 399486
rect 251088 399218 251130 399454
rect 251366 399218 251408 399454
rect 251088 399134 251408 399218
rect 251088 398898 251130 399134
rect 251366 398898 251408 399134
rect 251088 398866 251408 398898
rect 281808 399454 282128 399486
rect 281808 399218 281850 399454
rect 282086 399218 282128 399454
rect 281808 399134 282128 399218
rect 281808 398898 281850 399134
rect 282086 398898 282128 399134
rect 281808 398866 282128 398898
rect 312528 399454 312848 399486
rect 312528 399218 312570 399454
rect 312806 399218 312848 399454
rect 312528 399134 312848 399218
rect 312528 398898 312570 399134
rect 312806 398898 312848 399134
rect 312528 398866 312848 398898
rect 343248 399454 343568 399486
rect 343248 399218 343290 399454
rect 343526 399218 343568 399454
rect 343248 399134 343568 399218
rect 343248 398898 343290 399134
rect 343526 398898 343568 399134
rect 343248 398866 343568 398898
rect 373968 399454 374288 399486
rect 373968 399218 374010 399454
rect 374246 399218 374288 399454
rect 373968 399134 374288 399218
rect 373968 398898 374010 399134
rect 374246 398898 374288 399134
rect 373968 398866 374288 398898
rect 404688 399454 405008 399486
rect 404688 399218 404730 399454
rect 404966 399218 405008 399454
rect 404688 399134 405008 399218
rect 404688 398898 404730 399134
rect 404966 398898 405008 399134
rect 404688 398866 405008 398898
rect 435408 399454 435728 399486
rect 435408 399218 435450 399454
rect 435686 399218 435728 399454
rect 435408 399134 435728 399218
rect 435408 398898 435450 399134
rect 435686 398898 435728 399134
rect 435408 398866 435728 398898
rect 174288 381454 174608 381486
rect 174288 381218 174330 381454
rect 174566 381218 174608 381454
rect 174288 381134 174608 381218
rect 174288 380898 174330 381134
rect 174566 380898 174608 381134
rect 174288 380866 174608 380898
rect 205008 381454 205328 381486
rect 205008 381218 205050 381454
rect 205286 381218 205328 381454
rect 205008 381134 205328 381218
rect 205008 380898 205050 381134
rect 205286 380898 205328 381134
rect 205008 380866 205328 380898
rect 235728 381454 236048 381486
rect 235728 381218 235770 381454
rect 236006 381218 236048 381454
rect 235728 381134 236048 381218
rect 235728 380898 235770 381134
rect 236006 380898 236048 381134
rect 235728 380866 236048 380898
rect 266448 381454 266768 381486
rect 266448 381218 266490 381454
rect 266726 381218 266768 381454
rect 266448 381134 266768 381218
rect 266448 380898 266490 381134
rect 266726 380898 266768 381134
rect 266448 380866 266768 380898
rect 297168 381454 297488 381486
rect 297168 381218 297210 381454
rect 297446 381218 297488 381454
rect 297168 381134 297488 381218
rect 297168 380898 297210 381134
rect 297446 380898 297488 381134
rect 297168 380866 297488 380898
rect 327888 381454 328208 381486
rect 327888 381218 327930 381454
rect 328166 381218 328208 381454
rect 327888 381134 328208 381218
rect 327888 380898 327930 381134
rect 328166 380898 328208 381134
rect 327888 380866 328208 380898
rect 358608 381454 358928 381486
rect 358608 381218 358650 381454
rect 358886 381218 358928 381454
rect 358608 381134 358928 381218
rect 358608 380898 358650 381134
rect 358886 380898 358928 381134
rect 358608 380866 358928 380898
rect 389328 381454 389648 381486
rect 389328 381218 389370 381454
rect 389606 381218 389648 381454
rect 389328 381134 389648 381218
rect 389328 380898 389370 381134
rect 389606 380898 389648 381134
rect 389328 380866 389648 380898
rect 420048 381454 420368 381486
rect 420048 381218 420090 381454
rect 420326 381218 420368 381454
rect 420048 381134 420368 381218
rect 420048 380898 420090 381134
rect 420326 380898 420368 381134
rect 420048 380866 420368 380898
rect 158928 363454 159248 363486
rect 158928 363218 158970 363454
rect 159206 363218 159248 363454
rect 158928 363134 159248 363218
rect 158928 362898 158970 363134
rect 159206 362898 159248 363134
rect 158928 362866 159248 362898
rect 189648 363454 189968 363486
rect 189648 363218 189690 363454
rect 189926 363218 189968 363454
rect 189648 363134 189968 363218
rect 189648 362898 189690 363134
rect 189926 362898 189968 363134
rect 189648 362866 189968 362898
rect 220368 363454 220688 363486
rect 220368 363218 220410 363454
rect 220646 363218 220688 363454
rect 220368 363134 220688 363218
rect 220368 362898 220410 363134
rect 220646 362898 220688 363134
rect 220368 362866 220688 362898
rect 251088 363454 251408 363486
rect 251088 363218 251130 363454
rect 251366 363218 251408 363454
rect 251088 363134 251408 363218
rect 251088 362898 251130 363134
rect 251366 362898 251408 363134
rect 251088 362866 251408 362898
rect 281808 363454 282128 363486
rect 281808 363218 281850 363454
rect 282086 363218 282128 363454
rect 281808 363134 282128 363218
rect 281808 362898 281850 363134
rect 282086 362898 282128 363134
rect 281808 362866 282128 362898
rect 312528 363454 312848 363486
rect 312528 363218 312570 363454
rect 312806 363218 312848 363454
rect 312528 363134 312848 363218
rect 312528 362898 312570 363134
rect 312806 362898 312848 363134
rect 312528 362866 312848 362898
rect 343248 363454 343568 363486
rect 343248 363218 343290 363454
rect 343526 363218 343568 363454
rect 343248 363134 343568 363218
rect 343248 362898 343290 363134
rect 343526 362898 343568 363134
rect 343248 362866 343568 362898
rect 373968 363454 374288 363486
rect 373968 363218 374010 363454
rect 374246 363218 374288 363454
rect 373968 363134 374288 363218
rect 373968 362898 374010 363134
rect 374246 362898 374288 363134
rect 373968 362866 374288 362898
rect 404688 363454 405008 363486
rect 404688 363218 404730 363454
rect 404966 363218 405008 363454
rect 404688 363134 405008 363218
rect 404688 362898 404730 363134
rect 404966 362898 405008 363134
rect 404688 362866 405008 362898
rect 435408 363454 435728 363486
rect 435408 363218 435450 363454
rect 435686 363218 435728 363454
rect 435408 363134 435728 363218
rect 435408 362898 435450 363134
rect 435686 362898 435728 363134
rect 435408 362866 435728 362898
rect 174288 345454 174608 345486
rect 174288 345218 174330 345454
rect 174566 345218 174608 345454
rect 174288 345134 174608 345218
rect 174288 344898 174330 345134
rect 174566 344898 174608 345134
rect 174288 344866 174608 344898
rect 205008 345454 205328 345486
rect 205008 345218 205050 345454
rect 205286 345218 205328 345454
rect 205008 345134 205328 345218
rect 205008 344898 205050 345134
rect 205286 344898 205328 345134
rect 205008 344866 205328 344898
rect 235728 345454 236048 345486
rect 235728 345218 235770 345454
rect 236006 345218 236048 345454
rect 235728 345134 236048 345218
rect 235728 344898 235770 345134
rect 236006 344898 236048 345134
rect 235728 344866 236048 344898
rect 266448 345454 266768 345486
rect 266448 345218 266490 345454
rect 266726 345218 266768 345454
rect 266448 345134 266768 345218
rect 266448 344898 266490 345134
rect 266726 344898 266768 345134
rect 266448 344866 266768 344898
rect 297168 345454 297488 345486
rect 297168 345218 297210 345454
rect 297446 345218 297488 345454
rect 297168 345134 297488 345218
rect 297168 344898 297210 345134
rect 297446 344898 297488 345134
rect 297168 344866 297488 344898
rect 327888 345454 328208 345486
rect 327888 345218 327930 345454
rect 328166 345218 328208 345454
rect 327888 345134 328208 345218
rect 327888 344898 327930 345134
rect 328166 344898 328208 345134
rect 327888 344866 328208 344898
rect 358608 345454 358928 345486
rect 358608 345218 358650 345454
rect 358886 345218 358928 345454
rect 358608 345134 358928 345218
rect 358608 344898 358650 345134
rect 358886 344898 358928 345134
rect 358608 344866 358928 344898
rect 389328 345454 389648 345486
rect 389328 345218 389370 345454
rect 389606 345218 389648 345454
rect 389328 345134 389648 345218
rect 389328 344898 389370 345134
rect 389606 344898 389648 345134
rect 389328 344866 389648 344898
rect 420048 345454 420368 345486
rect 420048 345218 420090 345454
rect 420326 345218 420368 345454
rect 420048 345134 420368 345218
rect 420048 344898 420090 345134
rect 420326 344898 420368 345134
rect 420048 344866 420368 344898
rect 158928 327454 159248 327486
rect 158928 327218 158970 327454
rect 159206 327218 159248 327454
rect 158928 327134 159248 327218
rect 158928 326898 158970 327134
rect 159206 326898 159248 327134
rect 158928 326866 159248 326898
rect 189648 327454 189968 327486
rect 189648 327218 189690 327454
rect 189926 327218 189968 327454
rect 189648 327134 189968 327218
rect 189648 326898 189690 327134
rect 189926 326898 189968 327134
rect 189648 326866 189968 326898
rect 220368 327454 220688 327486
rect 220368 327218 220410 327454
rect 220646 327218 220688 327454
rect 220368 327134 220688 327218
rect 220368 326898 220410 327134
rect 220646 326898 220688 327134
rect 220368 326866 220688 326898
rect 251088 327454 251408 327486
rect 251088 327218 251130 327454
rect 251366 327218 251408 327454
rect 251088 327134 251408 327218
rect 251088 326898 251130 327134
rect 251366 326898 251408 327134
rect 251088 326866 251408 326898
rect 281808 327454 282128 327486
rect 281808 327218 281850 327454
rect 282086 327218 282128 327454
rect 281808 327134 282128 327218
rect 281808 326898 281850 327134
rect 282086 326898 282128 327134
rect 281808 326866 282128 326898
rect 312528 327454 312848 327486
rect 312528 327218 312570 327454
rect 312806 327218 312848 327454
rect 312528 327134 312848 327218
rect 312528 326898 312570 327134
rect 312806 326898 312848 327134
rect 312528 326866 312848 326898
rect 343248 327454 343568 327486
rect 343248 327218 343290 327454
rect 343526 327218 343568 327454
rect 343248 327134 343568 327218
rect 343248 326898 343290 327134
rect 343526 326898 343568 327134
rect 343248 326866 343568 326898
rect 373968 327454 374288 327486
rect 373968 327218 374010 327454
rect 374246 327218 374288 327454
rect 373968 327134 374288 327218
rect 373968 326898 374010 327134
rect 374246 326898 374288 327134
rect 373968 326866 374288 326898
rect 404688 327454 405008 327486
rect 404688 327218 404730 327454
rect 404966 327218 405008 327454
rect 404688 327134 405008 327218
rect 404688 326898 404730 327134
rect 404966 326898 405008 327134
rect 404688 326866 405008 326898
rect 435408 327454 435728 327486
rect 435408 327218 435450 327454
rect 435686 327218 435728 327454
rect 435408 327134 435728 327218
rect 435408 326898 435450 327134
rect 435686 326898 435728 327134
rect 435408 326866 435728 326898
rect 174288 309454 174608 309486
rect 174288 309218 174330 309454
rect 174566 309218 174608 309454
rect 174288 309134 174608 309218
rect 174288 308898 174330 309134
rect 174566 308898 174608 309134
rect 174288 308866 174608 308898
rect 205008 309454 205328 309486
rect 205008 309218 205050 309454
rect 205286 309218 205328 309454
rect 205008 309134 205328 309218
rect 205008 308898 205050 309134
rect 205286 308898 205328 309134
rect 205008 308866 205328 308898
rect 235728 309454 236048 309486
rect 235728 309218 235770 309454
rect 236006 309218 236048 309454
rect 235728 309134 236048 309218
rect 235728 308898 235770 309134
rect 236006 308898 236048 309134
rect 235728 308866 236048 308898
rect 266448 309454 266768 309486
rect 266448 309218 266490 309454
rect 266726 309218 266768 309454
rect 266448 309134 266768 309218
rect 266448 308898 266490 309134
rect 266726 308898 266768 309134
rect 266448 308866 266768 308898
rect 297168 309454 297488 309486
rect 297168 309218 297210 309454
rect 297446 309218 297488 309454
rect 297168 309134 297488 309218
rect 297168 308898 297210 309134
rect 297446 308898 297488 309134
rect 297168 308866 297488 308898
rect 327888 309454 328208 309486
rect 327888 309218 327930 309454
rect 328166 309218 328208 309454
rect 327888 309134 328208 309218
rect 327888 308898 327930 309134
rect 328166 308898 328208 309134
rect 327888 308866 328208 308898
rect 358608 309454 358928 309486
rect 358608 309218 358650 309454
rect 358886 309218 358928 309454
rect 358608 309134 358928 309218
rect 358608 308898 358650 309134
rect 358886 308898 358928 309134
rect 358608 308866 358928 308898
rect 389328 309454 389648 309486
rect 389328 309218 389370 309454
rect 389606 309218 389648 309454
rect 389328 309134 389648 309218
rect 389328 308898 389370 309134
rect 389606 308898 389648 309134
rect 389328 308866 389648 308898
rect 420048 309454 420368 309486
rect 420048 309218 420090 309454
rect 420326 309218 420368 309454
rect 420048 309134 420368 309218
rect 420048 308898 420090 309134
rect 420326 308898 420368 309134
rect 420048 308866 420368 308898
rect 158928 291454 159248 291486
rect 158928 291218 158970 291454
rect 159206 291218 159248 291454
rect 158928 291134 159248 291218
rect 158928 290898 158970 291134
rect 159206 290898 159248 291134
rect 158928 290866 159248 290898
rect 189648 291454 189968 291486
rect 189648 291218 189690 291454
rect 189926 291218 189968 291454
rect 189648 291134 189968 291218
rect 189648 290898 189690 291134
rect 189926 290898 189968 291134
rect 189648 290866 189968 290898
rect 220368 291454 220688 291486
rect 220368 291218 220410 291454
rect 220646 291218 220688 291454
rect 220368 291134 220688 291218
rect 220368 290898 220410 291134
rect 220646 290898 220688 291134
rect 220368 290866 220688 290898
rect 251088 291454 251408 291486
rect 251088 291218 251130 291454
rect 251366 291218 251408 291454
rect 251088 291134 251408 291218
rect 251088 290898 251130 291134
rect 251366 290898 251408 291134
rect 251088 290866 251408 290898
rect 281808 291454 282128 291486
rect 281808 291218 281850 291454
rect 282086 291218 282128 291454
rect 281808 291134 282128 291218
rect 281808 290898 281850 291134
rect 282086 290898 282128 291134
rect 281808 290866 282128 290898
rect 312528 291454 312848 291486
rect 312528 291218 312570 291454
rect 312806 291218 312848 291454
rect 312528 291134 312848 291218
rect 312528 290898 312570 291134
rect 312806 290898 312848 291134
rect 312528 290866 312848 290898
rect 343248 291454 343568 291486
rect 343248 291218 343290 291454
rect 343526 291218 343568 291454
rect 343248 291134 343568 291218
rect 343248 290898 343290 291134
rect 343526 290898 343568 291134
rect 343248 290866 343568 290898
rect 373968 291454 374288 291486
rect 373968 291218 374010 291454
rect 374246 291218 374288 291454
rect 373968 291134 374288 291218
rect 373968 290898 374010 291134
rect 374246 290898 374288 291134
rect 373968 290866 374288 290898
rect 404688 291454 405008 291486
rect 404688 291218 404730 291454
rect 404966 291218 405008 291454
rect 404688 291134 405008 291218
rect 404688 290898 404730 291134
rect 404966 290898 405008 291134
rect 404688 290866 405008 290898
rect 435408 291454 435728 291486
rect 435408 291218 435450 291454
rect 435686 291218 435728 291454
rect 435408 291134 435728 291218
rect 435408 290898 435450 291134
rect 435686 290898 435728 291134
rect 435408 290866 435728 290898
rect 174288 273454 174608 273486
rect 174288 273218 174330 273454
rect 174566 273218 174608 273454
rect 174288 273134 174608 273218
rect 174288 272898 174330 273134
rect 174566 272898 174608 273134
rect 174288 272866 174608 272898
rect 205008 273454 205328 273486
rect 205008 273218 205050 273454
rect 205286 273218 205328 273454
rect 205008 273134 205328 273218
rect 205008 272898 205050 273134
rect 205286 272898 205328 273134
rect 205008 272866 205328 272898
rect 235728 273454 236048 273486
rect 235728 273218 235770 273454
rect 236006 273218 236048 273454
rect 235728 273134 236048 273218
rect 235728 272898 235770 273134
rect 236006 272898 236048 273134
rect 235728 272866 236048 272898
rect 266448 273454 266768 273486
rect 266448 273218 266490 273454
rect 266726 273218 266768 273454
rect 266448 273134 266768 273218
rect 266448 272898 266490 273134
rect 266726 272898 266768 273134
rect 266448 272866 266768 272898
rect 297168 273454 297488 273486
rect 297168 273218 297210 273454
rect 297446 273218 297488 273454
rect 297168 273134 297488 273218
rect 297168 272898 297210 273134
rect 297446 272898 297488 273134
rect 297168 272866 297488 272898
rect 327888 273454 328208 273486
rect 327888 273218 327930 273454
rect 328166 273218 328208 273454
rect 327888 273134 328208 273218
rect 327888 272898 327930 273134
rect 328166 272898 328208 273134
rect 327888 272866 328208 272898
rect 358608 273454 358928 273486
rect 358608 273218 358650 273454
rect 358886 273218 358928 273454
rect 358608 273134 358928 273218
rect 358608 272898 358650 273134
rect 358886 272898 358928 273134
rect 358608 272866 358928 272898
rect 389328 273454 389648 273486
rect 389328 273218 389370 273454
rect 389606 273218 389648 273454
rect 389328 273134 389648 273218
rect 389328 272898 389370 273134
rect 389606 272898 389648 273134
rect 389328 272866 389648 272898
rect 420048 273454 420368 273486
rect 420048 273218 420090 273454
rect 420326 273218 420368 273454
rect 420048 273134 420368 273218
rect 420048 272898 420090 273134
rect 420326 272898 420368 273134
rect 420048 272866 420368 272898
rect 158928 255454 159248 255486
rect 158928 255218 158970 255454
rect 159206 255218 159248 255454
rect 158928 255134 159248 255218
rect 158928 254898 158970 255134
rect 159206 254898 159248 255134
rect 158928 254866 159248 254898
rect 189648 255454 189968 255486
rect 189648 255218 189690 255454
rect 189926 255218 189968 255454
rect 189648 255134 189968 255218
rect 189648 254898 189690 255134
rect 189926 254898 189968 255134
rect 189648 254866 189968 254898
rect 220368 255454 220688 255486
rect 220368 255218 220410 255454
rect 220646 255218 220688 255454
rect 220368 255134 220688 255218
rect 220368 254898 220410 255134
rect 220646 254898 220688 255134
rect 220368 254866 220688 254898
rect 251088 255454 251408 255486
rect 251088 255218 251130 255454
rect 251366 255218 251408 255454
rect 251088 255134 251408 255218
rect 251088 254898 251130 255134
rect 251366 254898 251408 255134
rect 251088 254866 251408 254898
rect 281808 255454 282128 255486
rect 281808 255218 281850 255454
rect 282086 255218 282128 255454
rect 281808 255134 282128 255218
rect 281808 254898 281850 255134
rect 282086 254898 282128 255134
rect 281808 254866 282128 254898
rect 312528 255454 312848 255486
rect 312528 255218 312570 255454
rect 312806 255218 312848 255454
rect 312528 255134 312848 255218
rect 312528 254898 312570 255134
rect 312806 254898 312848 255134
rect 312528 254866 312848 254898
rect 343248 255454 343568 255486
rect 343248 255218 343290 255454
rect 343526 255218 343568 255454
rect 343248 255134 343568 255218
rect 343248 254898 343290 255134
rect 343526 254898 343568 255134
rect 343248 254866 343568 254898
rect 373968 255454 374288 255486
rect 373968 255218 374010 255454
rect 374246 255218 374288 255454
rect 373968 255134 374288 255218
rect 373968 254898 374010 255134
rect 374246 254898 374288 255134
rect 373968 254866 374288 254898
rect 404688 255454 405008 255486
rect 404688 255218 404730 255454
rect 404966 255218 405008 255454
rect 404688 255134 405008 255218
rect 404688 254898 404730 255134
rect 404966 254898 405008 255134
rect 404688 254866 405008 254898
rect 435408 255454 435728 255486
rect 435408 255218 435450 255454
rect 435686 255218 435728 255454
rect 435408 255134 435728 255218
rect 435408 254898 435450 255134
rect 435686 254898 435728 255134
rect 435408 254866 435728 254898
rect 174288 237454 174608 237486
rect 174288 237218 174330 237454
rect 174566 237218 174608 237454
rect 174288 237134 174608 237218
rect 174288 236898 174330 237134
rect 174566 236898 174608 237134
rect 174288 236866 174608 236898
rect 205008 237454 205328 237486
rect 205008 237218 205050 237454
rect 205286 237218 205328 237454
rect 205008 237134 205328 237218
rect 205008 236898 205050 237134
rect 205286 236898 205328 237134
rect 205008 236866 205328 236898
rect 235728 237454 236048 237486
rect 235728 237218 235770 237454
rect 236006 237218 236048 237454
rect 235728 237134 236048 237218
rect 235728 236898 235770 237134
rect 236006 236898 236048 237134
rect 235728 236866 236048 236898
rect 266448 237454 266768 237486
rect 266448 237218 266490 237454
rect 266726 237218 266768 237454
rect 266448 237134 266768 237218
rect 266448 236898 266490 237134
rect 266726 236898 266768 237134
rect 266448 236866 266768 236898
rect 297168 237454 297488 237486
rect 297168 237218 297210 237454
rect 297446 237218 297488 237454
rect 297168 237134 297488 237218
rect 297168 236898 297210 237134
rect 297446 236898 297488 237134
rect 297168 236866 297488 236898
rect 327888 237454 328208 237486
rect 327888 237218 327930 237454
rect 328166 237218 328208 237454
rect 327888 237134 328208 237218
rect 327888 236898 327930 237134
rect 328166 236898 328208 237134
rect 327888 236866 328208 236898
rect 358608 237454 358928 237486
rect 358608 237218 358650 237454
rect 358886 237218 358928 237454
rect 358608 237134 358928 237218
rect 358608 236898 358650 237134
rect 358886 236898 358928 237134
rect 358608 236866 358928 236898
rect 389328 237454 389648 237486
rect 389328 237218 389370 237454
rect 389606 237218 389648 237454
rect 389328 237134 389648 237218
rect 389328 236898 389370 237134
rect 389606 236898 389648 237134
rect 389328 236866 389648 236898
rect 420048 237454 420368 237486
rect 420048 237218 420090 237454
rect 420326 237218 420368 237454
rect 420048 237134 420368 237218
rect 420048 236898 420090 237134
rect 420326 236898 420368 237134
rect 420048 236866 420368 236898
rect 158928 219454 159248 219486
rect 158928 219218 158970 219454
rect 159206 219218 159248 219454
rect 158928 219134 159248 219218
rect 158928 218898 158970 219134
rect 159206 218898 159248 219134
rect 158928 218866 159248 218898
rect 189648 219454 189968 219486
rect 189648 219218 189690 219454
rect 189926 219218 189968 219454
rect 189648 219134 189968 219218
rect 189648 218898 189690 219134
rect 189926 218898 189968 219134
rect 189648 218866 189968 218898
rect 220368 219454 220688 219486
rect 220368 219218 220410 219454
rect 220646 219218 220688 219454
rect 220368 219134 220688 219218
rect 220368 218898 220410 219134
rect 220646 218898 220688 219134
rect 220368 218866 220688 218898
rect 251088 219454 251408 219486
rect 251088 219218 251130 219454
rect 251366 219218 251408 219454
rect 251088 219134 251408 219218
rect 251088 218898 251130 219134
rect 251366 218898 251408 219134
rect 251088 218866 251408 218898
rect 281808 219454 282128 219486
rect 281808 219218 281850 219454
rect 282086 219218 282128 219454
rect 281808 219134 282128 219218
rect 281808 218898 281850 219134
rect 282086 218898 282128 219134
rect 281808 218866 282128 218898
rect 312528 219454 312848 219486
rect 312528 219218 312570 219454
rect 312806 219218 312848 219454
rect 312528 219134 312848 219218
rect 312528 218898 312570 219134
rect 312806 218898 312848 219134
rect 312528 218866 312848 218898
rect 343248 219454 343568 219486
rect 343248 219218 343290 219454
rect 343526 219218 343568 219454
rect 343248 219134 343568 219218
rect 343248 218898 343290 219134
rect 343526 218898 343568 219134
rect 343248 218866 343568 218898
rect 373968 219454 374288 219486
rect 373968 219218 374010 219454
rect 374246 219218 374288 219454
rect 373968 219134 374288 219218
rect 373968 218898 374010 219134
rect 374246 218898 374288 219134
rect 373968 218866 374288 218898
rect 404688 219454 405008 219486
rect 404688 219218 404730 219454
rect 404966 219218 405008 219454
rect 404688 219134 405008 219218
rect 404688 218898 404730 219134
rect 404966 218898 405008 219134
rect 404688 218866 405008 218898
rect 435408 219454 435728 219486
rect 435408 219218 435450 219454
rect 435686 219218 435728 219454
rect 435408 219134 435728 219218
rect 435408 218898 435450 219134
rect 435686 218898 435728 219134
rect 435408 218866 435728 218898
rect 174288 201454 174608 201486
rect 174288 201218 174330 201454
rect 174566 201218 174608 201454
rect 174288 201134 174608 201218
rect 174288 200898 174330 201134
rect 174566 200898 174608 201134
rect 174288 200866 174608 200898
rect 205008 201454 205328 201486
rect 205008 201218 205050 201454
rect 205286 201218 205328 201454
rect 205008 201134 205328 201218
rect 205008 200898 205050 201134
rect 205286 200898 205328 201134
rect 205008 200866 205328 200898
rect 235728 201454 236048 201486
rect 235728 201218 235770 201454
rect 236006 201218 236048 201454
rect 235728 201134 236048 201218
rect 235728 200898 235770 201134
rect 236006 200898 236048 201134
rect 235728 200866 236048 200898
rect 266448 201454 266768 201486
rect 266448 201218 266490 201454
rect 266726 201218 266768 201454
rect 266448 201134 266768 201218
rect 266448 200898 266490 201134
rect 266726 200898 266768 201134
rect 266448 200866 266768 200898
rect 297168 201454 297488 201486
rect 297168 201218 297210 201454
rect 297446 201218 297488 201454
rect 297168 201134 297488 201218
rect 297168 200898 297210 201134
rect 297446 200898 297488 201134
rect 297168 200866 297488 200898
rect 327888 201454 328208 201486
rect 327888 201218 327930 201454
rect 328166 201218 328208 201454
rect 327888 201134 328208 201218
rect 327888 200898 327930 201134
rect 328166 200898 328208 201134
rect 327888 200866 328208 200898
rect 358608 201454 358928 201486
rect 358608 201218 358650 201454
rect 358886 201218 358928 201454
rect 358608 201134 358928 201218
rect 358608 200898 358650 201134
rect 358886 200898 358928 201134
rect 358608 200866 358928 200898
rect 389328 201454 389648 201486
rect 389328 201218 389370 201454
rect 389606 201218 389648 201454
rect 389328 201134 389648 201218
rect 389328 200898 389370 201134
rect 389606 200898 389648 201134
rect 389328 200866 389648 200898
rect 420048 201454 420368 201486
rect 420048 201218 420090 201454
rect 420326 201218 420368 201454
rect 420048 201134 420368 201218
rect 420048 200898 420090 201134
rect 420326 200898 420368 201134
rect 420048 200866 420368 200898
rect 158928 183454 159248 183486
rect 158928 183218 158970 183454
rect 159206 183218 159248 183454
rect 158928 183134 159248 183218
rect 158928 182898 158970 183134
rect 159206 182898 159248 183134
rect 158928 182866 159248 182898
rect 189648 183454 189968 183486
rect 189648 183218 189690 183454
rect 189926 183218 189968 183454
rect 189648 183134 189968 183218
rect 189648 182898 189690 183134
rect 189926 182898 189968 183134
rect 189648 182866 189968 182898
rect 220368 183454 220688 183486
rect 220368 183218 220410 183454
rect 220646 183218 220688 183454
rect 220368 183134 220688 183218
rect 220368 182898 220410 183134
rect 220646 182898 220688 183134
rect 220368 182866 220688 182898
rect 251088 183454 251408 183486
rect 251088 183218 251130 183454
rect 251366 183218 251408 183454
rect 251088 183134 251408 183218
rect 251088 182898 251130 183134
rect 251366 182898 251408 183134
rect 251088 182866 251408 182898
rect 281808 183454 282128 183486
rect 281808 183218 281850 183454
rect 282086 183218 282128 183454
rect 281808 183134 282128 183218
rect 281808 182898 281850 183134
rect 282086 182898 282128 183134
rect 281808 182866 282128 182898
rect 312528 183454 312848 183486
rect 312528 183218 312570 183454
rect 312806 183218 312848 183454
rect 312528 183134 312848 183218
rect 312528 182898 312570 183134
rect 312806 182898 312848 183134
rect 312528 182866 312848 182898
rect 343248 183454 343568 183486
rect 343248 183218 343290 183454
rect 343526 183218 343568 183454
rect 343248 183134 343568 183218
rect 343248 182898 343290 183134
rect 343526 182898 343568 183134
rect 343248 182866 343568 182898
rect 373968 183454 374288 183486
rect 373968 183218 374010 183454
rect 374246 183218 374288 183454
rect 373968 183134 374288 183218
rect 373968 182898 374010 183134
rect 374246 182898 374288 183134
rect 373968 182866 374288 182898
rect 404688 183454 405008 183486
rect 404688 183218 404730 183454
rect 404966 183218 405008 183454
rect 404688 183134 405008 183218
rect 404688 182898 404730 183134
rect 404966 182898 405008 183134
rect 404688 182866 405008 182898
rect 435408 183454 435728 183486
rect 435408 183218 435450 183454
rect 435686 183218 435728 183454
rect 435408 183134 435728 183218
rect 435408 182898 435450 183134
rect 435686 182898 435728 183134
rect 435408 182866 435728 182898
rect 174288 165454 174608 165486
rect 174288 165218 174330 165454
rect 174566 165218 174608 165454
rect 174288 165134 174608 165218
rect 174288 164898 174330 165134
rect 174566 164898 174608 165134
rect 174288 164866 174608 164898
rect 205008 165454 205328 165486
rect 205008 165218 205050 165454
rect 205286 165218 205328 165454
rect 205008 165134 205328 165218
rect 205008 164898 205050 165134
rect 205286 164898 205328 165134
rect 205008 164866 205328 164898
rect 235728 165454 236048 165486
rect 235728 165218 235770 165454
rect 236006 165218 236048 165454
rect 235728 165134 236048 165218
rect 235728 164898 235770 165134
rect 236006 164898 236048 165134
rect 235728 164866 236048 164898
rect 266448 165454 266768 165486
rect 266448 165218 266490 165454
rect 266726 165218 266768 165454
rect 266448 165134 266768 165218
rect 266448 164898 266490 165134
rect 266726 164898 266768 165134
rect 266448 164866 266768 164898
rect 297168 165454 297488 165486
rect 297168 165218 297210 165454
rect 297446 165218 297488 165454
rect 297168 165134 297488 165218
rect 297168 164898 297210 165134
rect 297446 164898 297488 165134
rect 297168 164866 297488 164898
rect 327888 165454 328208 165486
rect 327888 165218 327930 165454
rect 328166 165218 328208 165454
rect 327888 165134 328208 165218
rect 327888 164898 327930 165134
rect 328166 164898 328208 165134
rect 327888 164866 328208 164898
rect 358608 165454 358928 165486
rect 358608 165218 358650 165454
rect 358886 165218 358928 165454
rect 358608 165134 358928 165218
rect 358608 164898 358650 165134
rect 358886 164898 358928 165134
rect 358608 164866 358928 164898
rect 389328 165454 389648 165486
rect 389328 165218 389370 165454
rect 389606 165218 389648 165454
rect 389328 165134 389648 165218
rect 389328 164898 389370 165134
rect 389606 164898 389648 165134
rect 389328 164866 389648 164898
rect 420048 165454 420368 165486
rect 420048 165218 420090 165454
rect 420326 165218 420368 165454
rect 420048 165134 420368 165218
rect 420048 164898 420090 165134
rect 420326 164898 420368 165134
rect 420048 164866 420368 164898
rect 158483 138140 158549 138141
rect 158483 138076 158484 138140
rect 158548 138076 158549 138140
rect 158483 138075 158549 138076
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 129454 164414 148400
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 133174 168134 148400
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 136894 171854 148400
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 140614 175574 148400
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 147454 182414 148400
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 115174 186134 148400
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 118894 189854 148400
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 122614 193574 148400
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 129454 200414 148400
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 133174 204134 148400
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 136894 207854 148400
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 140614 211574 148400
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 147454 218414 148400
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 115174 222134 148400
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 118894 225854 148400
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 122614 229574 148400
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 129454 236414 148400
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 133174 240134 148400
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 136894 243854 148400
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 140614 247574 148400
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 147454 254414 148400
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 115174 258134 148400
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 118894 261854 148400
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 122614 265574 148400
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 129454 272414 148400
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 133174 276134 148400
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 136894 279854 148400
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 140614 283574 148400
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 147454 290414 148400
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 115174 294134 148400
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 118894 297854 148400
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 122614 301574 148400
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 129454 308414 148400
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 133174 312134 148400
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 136894 315854 148400
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 140614 319574 148400
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 147454 326414 148400
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 115174 330134 148400
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 118894 333854 148400
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 122614 337574 148400
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 129454 344414 148400
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 133174 348134 148400
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 136894 351854 148400
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 140614 355574 148400
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 147454 362414 148400
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 115174 366134 148400
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 118894 369854 148400
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 122614 373574 148400
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 129454 380414 148400
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 133174 384134 148400
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 136894 387854 148400
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 140614 391574 148400
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 147454 398414 148400
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 115174 402134 148400
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 118894 405854 148400
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 122614 409574 148400
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 129454 416414 148400
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 133174 420134 148400
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 136894 423854 148400
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 140614 427574 148400
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 147454 434414 148400
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 436142 111757 436202 557499
rect 437514 115174 438134 148400
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 436139 111756 436205 111757
rect 436139 111692 436140 111756
rect 436204 111692 436205 111756
rect 436139 111691 436205 111692
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 79174 438134 114618
rect 438902 85509 438962 557499
rect 441234 118894 441854 148400
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 438899 85508 438965 85509
rect 438899 85444 438900 85508
rect 438964 85444 438965 85508
rect 438899 85443 438965 85444
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 82894 441854 118338
rect 442950 97885 443010 557499
rect 444954 122614 445574 148400
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 442947 97884 443013 97885
rect 442947 97820 442948 97884
rect 443012 97820 443013 97884
rect 442947 97819 443013 97820
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 445710 71773 445770 557499
rect 445707 71772 445773 71773
rect 445707 71708 445708 71772
rect 445772 71708 445773 71772
rect 445707 71707 445773 71708
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 448470 45525 448530 557499
rect 451046 557490 451290 557499
rect 451046 555930 451106 557490
rect 451046 555870 451474 555930
rect 450768 525454 451088 525486
rect 450768 525218 450810 525454
rect 451046 525218 451088 525454
rect 450768 525134 451088 525218
rect 450768 524898 450810 525134
rect 451046 524898 451088 525134
rect 450768 524866 451088 524898
rect 450768 489454 451088 489486
rect 450768 489218 450810 489454
rect 451046 489218 451088 489454
rect 450768 489134 451088 489218
rect 450768 488898 450810 489134
rect 451046 488898 451088 489134
rect 450768 488866 451088 488898
rect 450768 453454 451088 453486
rect 450768 453218 450810 453454
rect 451046 453218 451088 453454
rect 450768 453134 451088 453218
rect 450768 452898 450810 453134
rect 451046 452898 451088 453134
rect 450768 452866 451088 452898
rect 450768 417454 451088 417486
rect 450768 417218 450810 417454
rect 451046 417218 451088 417454
rect 450768 417134 451088 417218
rect 450768 416898 450810 417134
rect 451046 416898 451088 417134
rect 450768 416866 451088 416898
rect 450768 381454 451088 381486
rect 450768 381218 450810 381454
rect 451046 381218 451088 381454
rect 450768 381134 451088 381218
rect 450768 380898 450810 381134
rect 451046 380898 451088 381134
rect 450768 380866 451088 380898
rect 450768 345454 451088 345486
rect 450768 345218 450810 345454
rect 451046 345218 451088 345454
rect 450768 345134 451088 345218
rect 450768 344898 450810 345134
rect 451046 344898 451088 345134
rect 450768 344866 451088 344898
rect 450768 309454 451088 309486
rect 450768 309218 450810 309454
rect 451046 309218 451088 309454
rect 450768 309134 451088 309218
rect 450768 308898 450810 309134
rect 451046 308898 451088 309134
rect 450768 308866 451088 308898
rect 450768 273454 451088 273486
rect 450768 273218 450810 273454
rect 451046 273218 451088 273454
rect 450768 273134 451088 273218
rect 450768 272898 450810 273134
rect 451046 272898 451088 273134
rect 450768 272866 451088 272898
rect 450768 237454 451088 237486
rect 450768 237218 450810 237454
rect 451046 237218 451088 237454
rect 450768 237134 451088 237218
rect 450768 236898 450810 237134
rect 451046 236898 451088 237134
rect 450768 236866 451088 236898
rect 450768 201454 451088 201486
rect 450768 201218 450810 201454
rect 451046 201218 451088 201454
rect 450768 201134 451088 201218
rect 450768 200898 450810 201134
rect 451046 200898 451088 201134
rect 450768 200866 451088 200898
rect 450768 165454 451088 165486
rect 450768 165218 450810 165454
rect 451046 165218 451088 165454
rect 450768 165134 451088 165218
rect 450768 164898 450810 165134
rect 451046 164898 451088 165134
rect 450768 164866 451088 164898
rect 451414 151830 451474 555870
rect 451046 151770 451474 151830
rect 451046 59261 451106 151770
rect 451794 129454 452414 148400
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451043 59260 451109 59261
rect 451043 59196 451044 59260
rect 451108 59196 451109 59260
rect 451043 59195 451109 59196
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 448467 45524 448533 45525
rect 448467 45460 448468 45524
rect 448532 45460 448533 45524
rect 448467 45459 448533 45460
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 21454 452414 56898
rect 454174 33149 454234 557499
rect 455514 133174 456134 148400
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 454171 33148 454237 33149
rect 454171 33084 454172 33148
rect 454236 33084 454237 33148
rect 454171 33083 454237 33084
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 456750 6901 456810 557499
rect 459234 136894 459854 148400
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 456747 6900 456813 6901
rect 456747 6836 456748 6900
rect 456812 6836 456813 6900
rect 456747 6835 456813 6836
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 -5146 459854 28338
rect 460062 20637 460122 557499
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 462954 140614 463574 148400
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 460059 20636 460125 20637
rect 460059 20572 460060 20636
rect 460124 20572 460125 20636
rect 460059 20571 460125 20572
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 128250 543218 128486 543454
rect 128250 542898 128486 543134
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 128250 507218 128486 507454
rect 128250 506898 128486 507134
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 128250 471218 128486 471454
rect 128250 470898 128486 471134
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 128250 435218 128486 435454
rect 128250 434898 128486 435134
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 128250 399218 128486 399454
rect 128250 398898 128486 399134
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 128250 363218 128486 363454
rect 128250 362898 128486 363134
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 128250 327218 128486 327454
rect 128250 326898 128486 327134
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 128250 291218 128486 291454
rect 128250 290898 128486 291134
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 128250 255218 128486 255454
rect 128250 254898 128486 255134
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 128250 219218 128486 219454
rect 128250 218898 128486 219134
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 128250 183218 128486 183454
rect 128250 182898 128486 183134
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 143610 525218 143846 525454
rect 143610 524898 143846 525134
rect 143610 489218 143846 489454
rect 143610 488898 143846 489134
rect 143610 453218 143846 453454
rect 143610 452898 143846 453134
rect 143610 417218 143846 417454
rect 143610 416898 143846 417134
rect 143610 381218 143846 381454
rect 143610 380898 143846 381134
rect 143610 345218 143846 345454
rect 143610 344898 143846 345134
rect 143610 309218 143846 309454
rect 143610 308898 143846 309134
rect 143610 273218 143846 273454
rect 143610 272898 143846 273134
rect 143610 237218 143846 237454
rect 143610 236898 143846 237134
rect 143610 201218 143846 201454
rect 143610 200898 143846 201134
rect 143610 165218 143846 165454
rect 143610 164898 143846 165134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 158970 543218 159206 543454
rect 158970 542898 159206 543134
rect 189690 543218 189926 543454
rect 189690 542898 189926 543134
rect 220410 543218 220646 543454
rect 220410 542898 220646 543134
rect 251130 543218 251366 543454
rect 251130 542898 251366 543134
rect 281850 543218 282086 543454
rect 281850 542898 282086 543134
rect 312570 543218 312806 543454
rect 312570 542898 312806 543134
rect 343290 543218 343526 543454
rect 343290 542898 343526 543134
rect 374010 543218 374246 543454
rect 374010 542898 374246 543134
rect 404730 543218 404966 543454
rect 404730 542898 404966 543134
rect 435450 543218 435686 543454
rect 435450 542898 435686 543134
rect 174330 525218 174566 525454
rect 174330 524898 174566 525134
rect 205050 525218 205286 525454
rect 205050 524898 205286 525134
rect 235770 525218 236006 525454
rect 235770 524898 236006 525134
rect 266490 525218 266726 525454
rect 266490 524898 266726 525134
rect 297210 525218 297446 525454
rect 297210 524898 297446 525134
rect 327930 525218 328166 525454
rect 327930 524898 328166 525134
rect 358650 525218 358886 525454
rect 358650 524898 358886 525134
rect 389370 525218 389606 525454
rect 389370 524898 389606 525134
rect 420090 525218 420326 525454
rect 420090 524898 420326 525134
rect 158970 507218 159206 507454
rect 158970 506898 159206 507134
rect 189690 507218 189926 507454
rect 189690 506898 189926 507134
rect 220410 507218 220646 507454
rect 220410 506898 220646 507134
rect 251130 507218 251366 507454
rect 251130 506898 251366 507134
rect 281850 507218 282086 507454
rect 281850 506898 282086 507134
rect 312570 507218 312806 507454
rect 312570 506898 312806 507134
rect 343290 507218 343526 507454
rect 343290 506898 343526 507134
rect 374010 507218 374246 507454
rect 374010 506898 374246 507134
rect 404730 507218 404966 507454
rect 404730 506898 404966 507134
rect 435450 507218 435686 507454
rect 435450 506898 435686 507134
rect 174330 489218 174566 489454
rect 174330 488898 174566 489134
rect 205050 489218 205286 489454
rect 205050 488898 205286 489134
rect 235770 489218 236006 489454
rect 235770 488898 236006 489134
rect 266490 489218 266726 489454
rect 266490 488898 266726 489134
rect 297210 489218 297446 489454
rect 297210 488898 297446 489134
rect 327930 489218 328166 489454
rect 327930 488898 328166 489134
rect 358650 489218 358886 489454
rect 358650 488898 358886 489134
rect 389370 489218 389606 489454
rect 389370 488898 389606 489134
rect 420090 489218 420326 489454
rect 420090 488898 420326 489134
rect 158970 471218 159206 471454
rect 158970 470898 159206 471134
rect 189690 471218 189926 471454
rect 189690 470898 189926 471134
rect 220410 471218 220646 471454
rect 220410 470898 220646 471134
rect 251130 471218 251366 471454
rect 251130 470898 251366 471134
rect 281850 471218 282086 471454
rect 281850 470898 282086 471134
rect 312570 471218 312806 471454
rect 312570 470898 312806 471134
rect 343290 471218 343526 471454
rect 343290 470898 343526 471134
rect 374010 471218 374246 471454
rect 374010 470898 374246 471134
rect 404730 471218 404966 471454
rect 404730 470898 404966 471134
rect 435450 471218 435686 471454
rect 435450 470898 435686 471134
rect 174330 453218 174566 453454
rect 174330 452898 174566 453134
rect 205050 453218 205286 453454
rect 205050 452898 205286 453134
rect 235770 453218 236006 453454
rect 235770 452898 236006 453134
rect 266490 453218 266726 453454
rect 266490 452898 266726 453134
rect 297210 453218 297446 453454
rect 297210 452898 297446 453134
rect 327930 453218 328166 453454
rect 327930 452898 328166 453134
rect 358650 453218 358886 453454
rect 358650 452898 358886 453134
rect 389370 453218 389606 453454
rect 389370 452898 389606 453134
rect 420090 453218 420326 453454
rect 420090 452898 420326 453134
rect 158970 435218 159206 435454
rect 158970 434898 159206 435134
rect 189690 435218 189926 435454
rect 189690 434898 189926 435134
rect 220410 435218 220646 435454
rect 220410 434898 220646 435134
rect 251130 435218 251366 435454
rect 251130 434898 251366 435134
rect 281850 435218 282086 435454
rect 281850 434898 282086 435134
rect 312570 435218 312806 435454
rect 312570 434898 312806 435134
rect 343290 435218 343526 435454
rect 343290 434898 343526 435134
rect 374010 435218 374246 435454
rect 374010 434898 374246 435134
rect 404730 435218 404966 435454
rect 404730 434898 404966 435134
rect 435450 435218 435686 435454
rect 435450 434898 435686 435134
rect 174330 417218 174566 417454
rect 174330 416898 174566 417134
rect 205050 417218 205286 417454
rect 205050 416898 205286 417134
rect 235770 417218 236006 417454
rect 235770 416898 236006 417134
rect 266490 417218 266726 417454
rect 266490 416898 266726 417134
rect 297210 417218 297446 417454
rect 297210 416898 297446 417134
rect 327930 417218 328166 417454
rect 327930 416898 328166 417134
rect 358650 417218 358886 417454
rect 358650 416898 358886 417134
rect 389370 417218 389606 417454
rect 389370 416898 389606 417134
rect 420090 417218 420326 417454
rect 420090 416898 420326 417134
rect 158970 399218 159206 399454
rect 158970 398898 159206 399134
rect 189690 399218 189926 399454
rect 189690 398898 189926 399134
rect 220410 399218 220646 399454
rect 220410 398898 220646 399134
rect 251130 399218 251366 399454
rect 251130 398898 251366 399134
rect 281850 399218 282086 399454
rect 281850 398898 282086 399134
rect 312570 399218 312806 399454
rect 312570 398898 312806 399134
rect 343290 399218 343526 399454
rect 343290 398898 343526 399134
rect 374010 399218 374246 399454
rect 374010 398898 374246 399134
rect 404730 399218 404966 399454
rect 404730 398898 404966 399134
rect 435450 399218 435686 399454
rect 435450 398898 435686 399134
rect 174330 381218 174566 381454
rect 174330 380898 174566 381134
rect 205050 381218 205286 381454
rect 205050 380898 205286 381134
rect 235770 381218 236006 381454
rect 235770 380898 236006 381134
rect 266490 381218 266726 381454
rect 266490 380898 266726 381134
rect 297210 381218 297446 381454
rect 297210 380898 297446 381134
rect 327930 381218 328166 381454
rect 327930 380898 328166 381134
rect 358650 381218 358886 381454
rect 358650 380898 358886 381134
rect 389370 381218 389606 381454
rect 389370 380898 389606 381134
rect 420090 381218 420326 381454
rect 420090 380898 420326 381134
rect 158970 363218 159206 363454
rect 158970 362898 159206 363134
rect 189690 363218 189926 363454
rect 189690 362898 189926 363134
rect 220410 363218 220646 363454
rect 220410 362898 220646 363134
rect 251130 363218 251366 363454
rect 251130 362898 251366 363134
rect 281850 363218 282086 363454
rect 281850 362898 282086 363134
rect 312570 363218 312806 363454
rect 312570 362898 312806 363134
rect 343290 363218 343526 363454
rect 343290 362898 343526 363134
rect 374010 363218 374246 363454
rect 374010 362898 374246 363134
rect 404730 363218 404966 363454
rect 404730 362898 404966 363134
rect 435450 363218 435686 363454
rect 435450 362898 435686 363134
rect 174330 345218 174566 345454
rect 174330 344898 174566 345134
rect 205050 345218 205286 345454
rect 205050 344898 205286 345134
rect 235770 345218 236006 345454
rect 235770 344898 236006 345134
rect 266490 345218 266726 345454
rect 266490 344898 266726 345134
rect 297210 345218 297446 345454
rect 297210 344898 297446 345134
rect 327930 345218 328166 345454
rect 327930 344898 328166 345134
rect 358650 345218 358886 345454
rect 358650 344898 358886 345134
rect 389370 345218 389606 345454
rect 389370 344898 389606 345134
rect 420090 345218 420326 345454
rect 420090 344898 420326 345134
rect 158970 327218 159206 327454
rect 158970 326898 159206 327134
rect 189690 327218 189926 327454
rect 189690 326898 189926 327134
rect 220410 327218 220646 327454
rect 220410 326898 220646 327134
rect 251130 327218 251366 327454
rect 251130 326898 251366 327134
rect 281850 327218 282086 327454
rect 281850 326898 282086 327134
rect 312570 327218 312806 327454
rect 312570 326898 312806 327134
rect 343290 327218 343526 327454
rect 343290 326898 343526 327134
rect 374010 327218 374246 327454
rect 374010 326898 374246 327134
rect 404730 327218 404966 327454
rect 404730 326898 404966 327134
rect 435450 327218 435686 327454
rect 435450 326898 435686 327134
rect 174330 309218 174566 309454
rect 174330 308898 174566 309134
rect 205050 309218 205286 309454
rect 205050 308898 205286 309134
rect 235770 309218 236006 309454
rect 235770 308898 236006 309134
rect 266490 309218 266726 309454
rect 266490 308898 266726 309134
rect 297210 309218 297446 309454
rect 297210 308898 297446 309134
rect 327930 309218 328166 309454
rect 327930 308898 328166 309134
rect 358650 309218 358886 309454
rect 358650 308898 358886 309134
rect 389370 309218 389606 309454
rect 389370 308898 389606 309134
rect 420090 309218 420326 309454
rect 420090 308898 420326 309134
rect 158970 291218 159206 291454
rect 158970 290898 159206 291134
rect 189690 291218 189926 291454
rect 189690 290898 189926 291134
rect 220410 291218 220646 291454
rect 220410 290898 220646 291134
rect 251130 291218 251366 291454
rect 251130 290898 251366 291134
rect 281850 291218 282086 291454
rect 281850 290898 282086 291134
rect 312570 291218 312806 291454
rect 312570 290898 312806 291134
rect 343290 291218 343526 291454
rect 343290 290898 343526 291134
rect 374010 291218 374246 291454
rect 374010 290898 374246 291134
rect 404730 291218 404966 291454
rect 404730 290898 404966 291134
rect 435450 291218 435686 291454
rect 435450 290898 435686 291134
rect 174330 273218 174566 273454
rect 174330 272898 174566 273134
rect 205050 273218 205286 273454
rect 205050 272898 205286 273134
rect 235770 273218 236006 273454
rect 235770 272898 236006 273134
rect 266490 273218 266726 273454
rect 266490 272898 266726 273134
rect 297210 273218 297446 273454
rect 297210 272898 297446 273134
rect 327930 273218 328166 273454
rect 327930 272898 328166 273134
rect 358650 273218 358886 273454
rect 358650 272898 358886 273134
rect 389370 273218 389606 273454
rect 389370 272898 389606 273134
rect 420090 273218 420326 273454
rect 420090 272898 420326 273134
rect 158970 255218 159206 255454
rect 158970 254898 159206 255134
rect 189690 255218 189926 255454
rect 189690 254898 189926 255134
rect 220410 255218 220646 255454
rect 220410 254898 220646 255134
rect 251130 255218 251366 255454
rect 251130 254898 251366 255134
rect 281850 255218 282086 255454
rect 281850 254898 282086 255134
rect 312570 255218 312806 255454
rect 312570 254898 312806 255134
rect 343290 255218 343526 255454
rect 343290 254898 343526 255134
rect 374010 255218 374246 255454
rect 374010 254898 374246 255134
rect 404730 255218 404966 255454
rect 404730 254898 404966 255134
rect 435450 255218 435686 255454
rect 435450 254898 435686 255134
rect 174330 237218 174566 237454
rect 174330 236898 174566 237134
rect 205050 237218 205286 237454
rect 205050 236898 205286 237134
rect 235770 237218 236006 237454
rect 235770 236898 236006 237134
rect 266490 237218 266726 237454
rect 266490 236898 266726 237134
rect 297210 237218 297446 237454
rect 297210 236898 297446 237134
rect 327930 237218 328166 237454
rect 327930 236898 328166 237134
rect 358650 237218 358886 237454
rect 358650 236898 358886 237134
rect 389370 237218 389606 237454
rect 389370 236898 389606 237134
rect 420090 237218 420326 237454
rect 420090 236898 420326 237134
rect 158970 219218 159206 219454
rect 158970 218898 159206 219134
rect 189690 219218 189926 219454
rect 189690 218898 189926 219134
rect 220410 219218 220646 219454
rect 220410 218898 220646 219134
rect 251130 219218 251366 219454
rect 251130 218898 251366 219134
rect 281850 219218 282086 219454
rect 281850 218898 282086 219134
rect 312570 219218 312806 219454
rect 312570 218898 312806 219134
rect 343290 219218 343526 219454
rect 343290 218898 343526 219134
rect 374010 219218 374246 219454
rect 374010 218898 374246 219134
rect 404730 219218 404966 219454
rect 404730 218898 404966 219134
rect 435450 219218 435686 219454
rect 435450 218898 435686 219134
rect 174330 201218 174566 201454
rect 174330 200898 174566 201134
rect 205050 201218 205286 201454
rect 205050 200898 205286 201134
rect 235770 201218 236006 201454
rect 235770 200898 236006 201134
rect 266490 201218 266726 201454
rect 266490 200898 266726 201134
rect 297210 201218 297446 201454
rect 297210 200898 297446 201134
rect 327930 201218 328166 201454
rect 327930 200898 328166 201134
rect 358650 201218 358886 201454
rect 358650 200898 358886 201134
rect 389370 201218 389606 201454
rect 389370 200898 389606 201134
rect 420090 201218 420326 201454
rect 420090 200898 420326 201134
rect 158970 183218 159206 183454
rect 158970 182898 159206 183134
rect 189690 183218 189926 183454
rect 189690 182898 189926 183134
rect 220410 183218 220646 183454
rect 220410 182898 220646 183134
rect 251130 183218 251366 183454
rect 251130 182898 251366 183134
rect 281850 183218 282086 183454
rect 281850 182898 282086 183134
rect 312570 183218 312806 183454
rect 312570 182898 312806 183134
rect 343290 183218 343526 183454
rect 343290 182898 343526 183134
rect 374010 183218 374246 183454
rect 374010 182898 374246 183134
rect 404730 183218 404966 183454
rect 404730 182898 404966 183134
rect 435450 183218 435686 183454
rect 435450 182898 435686 183134
rect 174330 165218 174566 165454
rect 174330 164898 174566 165134
rect 205050 165218 205286 165454
rect 205050 164898 205286 165134
rect 235770 165218 236006 165454
rect 235770 164898 236006 165134
rect 266490 165218 266726 165454
rect 266490 164898 266726 165134
rect 297210 165218 297446 165454
rect 297210 164898 297446 165134
rect 327930 165218 328166 165454
rect 327930 164898 328166 165134
rect 358650 165218 358886 165454
rect 358650 164898 358886 165134
rect 389370 165218 389606 165454
rect 389370 164898 389606 165134
rect 420090 165218 420326 165454
rect 420090 164898 420326 165134
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 450810 525218 451046 525454
rect 450810 524898 451046 525134
rect 450810 489218 451046 489454
rect 450810 488898 451046 489134
rect 450810 453218 451046 453454
rect 450810 452898 451046 453134
rect 450810 417218 451046 417454
rect 450810 416898 451046 417134
rect 450810 381218 451046 381454
rect 450810 380898 451046 381134
rect 450810 345218 451046 345454
rect 450810 344898 451046 345134
rect 450810 309218 451046 309454
rect 450810 308898 451046 309134
rect 450810 273218 451046 273454
rect 450810 272898 451046 273134
rect 450810 237218 451046 237454
rect 450810 236898 451046 237134
rect 450810 201218 451046 201454
rect 450810 200898 451046 201134
rect 450810 165218 451046 165454
rect 450810 164898 451046 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 128250 543454
rect 128486 543218 158970 543454
rect 159206 543218 189690 543454
rect 189926 543218 220410 543454
rect 220646 543218 251130 543454
rect 251366 543218 281850 543454
rect 282086 543218 312570 543454
rect 312806 543218 343290 543454
rect 343526 543218 374010 543454
rect 374246 543218 404730 543454
rect 404966 543218 435450 543454
rect 435686 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 128250 543134
rect 128486 542898 158970 543134
rect 159206 542898 189690 543134
rect 189926 542898 220410 543134
rect 220646 542898 251130 543134
rect 251366 542898 281850 543134
rect 282086 542898 312570 543134
rect 312806 542898 343290 543134
rect 343526 542898 374010 543134
rect 374246 542898 404730 543134
rect 404966 542898 435450 543134
rect 435686 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 143610 525454
rect 143846 525218 174330 525454
rect 174566 525218 205050 525454
rect 205286 525218 235770 525454
rect 236006 525218 266490 525454
rect 266726 525218 297210 525454
rect 297446 525218 327930 525454
rect 328166 525218 358650 525454
rect 358886 525218 389370 525454
rect 389606 525218 420090 525454
rect 420326 525218 450810 525454
rect 451046 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 143610 525134
rect 143846 524898 174330 525134
rect 174566 524898 205050 525134
rect 205286 524898 235770 525134
rect 236006 524898 266490 525134
rect 266726 524898 297210 525134
rect 297446 524898 327930 525134
rect 328166 524898 358650 525134
rect 358886 524898 389370 525134
rect 389606 524898 420090 525134
rect 420326 524898 450810 525134
rect 451046 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 128250 507454
rect 128486 507218 158970 507454
rect 159206 507218 189690 507454
rect 189926 507218 220410 507454
rect 220646 507218 251130 507454
rect 251366 507218 281850 507454
rect 282086 507218 312570 507454
rect 312806 507218 343290 507454
rect 343526 507218 374010 507454
rect 374246 507218 404730 507454
rect 404966 507218 435450 507454
rect 435686 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 128250 507134
rect 128486 506898 158970 507134
rect 159206 506898 189690 507134
rect 189926 506898 220410 507134
rect 220646 506898 251130 507134
rect 251366 506898 281850 507134
rect 282086 506898 312570 507134
rect 312806 506898 343290 507134
rect 343526 506898 374010 507134
rect 374246 506898 404730 507134
rect 404966 506898 435450 507134
rect 435686 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 143610 489454
rect 143846 489218 174330 489454
rect 174566 489218 205050 489454
rect 205286 489218 235770 489454
rect 236006 489218 266490 489454
rect 266726 489218 297210 489454
rect 297446 489218 327930 489454
rect 328166 489218 358650 489454
rect 358886 489218 389370 489454
rect 389606 489218 420090 489454
rect 420326 489218 450810 489454
rect 451046 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 143610 489134
rect 143846 488898 174330 489134
rect 174566 488898 205050 489134
rect 205286 488898 235770 489134
rect 236006 488898 266490 489134
rect 266726 488898 297210 489134
rect 297446 488898 327930 489134
rect 328166 488898 358650 489134
rect 358886 488898 389370 489134
rect 389606 488898 420090 489134
rect 420326 488898 450810 489134
rect 451046 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 128250 471454
rect 128486 471218 158970 471454
rect 159206 471218 189690 471454
rect 189926 471218 220410 471454
rect 220646 471218 251130 471454
rect 251366 471218 281850 471454
rect 282086 471218 312570 471454
rect 312806 471218 343290 471454
rect 343526 471218 374010 471454
rect 374246 471218 404730 471454
rect 404966 471218 435450 471454
rect 435686 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 128250 471134
rect 128486 470898 158970 471134
rect 159206 470898 189690 471134
rect 189926 470898 220410 471134
rect 220646 470898 251130 471134
rect 251366 470898 281850 471134
rect 282086 470898 312570 471134
rect 312806 470898 343290 471134
rect 343526 470898 374010 471134
rect 374246 470898 404730 471134
rect 404966 470898 435450 471134
rect 435686 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 143610 453454
rect 143846 453218 174330 453454
rect 174566 453218 205050 453454
rect 205286 453218 235770 453454
rect 236006 453218 266490 453454
rect 266726 453218 297210 453454
rect 297446 453218 327930 453454
rect 328166 453218 358650 453454
rect 358886 453218 389370 453454
rect 389606 453218 420090 453454
rect 420326 453218 450810 453454
rect 451046 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 143610 453134
rect 143846 452898 174330 453134
rect 174566 452898 205050 453134
rect 205286 452898 235770 453134
rect 236006 452898 266490 453134
rect 266726 452898 297210 453134
rect 297446 452898 327930 453134
rect 328166 452898 358650 453134
rect 358886 452898 389370 453134
rect 389606 452898 420090 453134
rect 420326 452898 450810 453134
rect 451046 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 128250 435454
rect 128486 435218 158970 435454
rect 159206 435218 189690 435454
rect 189926 435218 220410 435454
rect 220646 435218 251130 435454
rect 251366 435218 281850 435454
rect 282086 435218 312570 435454
rect 312806 435218 343290 435454
rect 343526 435218 374010 435454
rect 374246 435218 404730 435454
rect 404966 435218 435450 435454
rect 435686 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 128250 435134
rect 128486 434898 158970 435134
rect 159206 434898 189690 435134
rect 189926 434898 220410 435134
rect 220646 434898 251130 435134
rect 251366 434898 281850 435134
rect 282086 434898 312570 435134
rect 312806 434898 343290 435134
rect 343526 434898 374010 435134
rect 374246 434898 404730 435134
rect 404966 434898 435450 435134
rect 435686 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 143610 417454
rect 143846 417218 174330 417454
rect 174566 417218 205050 417454
rect 205286 417218 235770 417454
rect 236006 417218 266490 417454
rect 266726 417218 297210 417454
rect 297446 417218 327930 417454
rect 328166 417218 358650 417454
rect 358886 417218 389370 417454
rect 389606 417218 420090 417454
rect 420326 417218 450810 417454
rect 451046 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 143610 417134
rect 143846 416898 174330 417134
rect 174566 416898 205050 417134
rect 205286 416898 235770 417134
rect 236006 416898 266490 417134
rect 266726 416898 297210 417134
rect 297446 416898 327930 417134
rect 328166 416898 358650 417134
rect 358886 416898 389370 417134
rect 389606 416898 420090 417134
rect 420326 416898 450810 417134
rect 451046 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 128250 399454
rect 128486 399218 158970 399454
rect 159206 399218 189690 399454
rect 189926 399218 220410 399454
rect 220646 399218 251130 399454
rect 251366 399218 281850 399454
rect 282086 399218 312570 399454
rect 312806 399218 343290 399454
rect 343526 399218 374010 399454
rect 374246 399218 404730 399454
rect 404966 399218 435450 399454
rect 435686 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 128250 399134
rect 128486 398898 158970 399134
rect 159206 398898 189690 399134
rect 189926 398898 220410 399134
rect 220646 398898 251130 399134
rect 251366 398898 281850 399134
rect 282086 398898 312570 399134
rect 312806 398898 343290 399134
rect 343526 398898 374010 399134
rect 374246 398898 404730 399134
rect 404966 398898 435450 399134
rect 435686 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 143610 381454
rect 143846 381218 174330 381454
rect 174566 381218 205050 381454
rect 205286 381218 235770 381454
rect 236006 381218 266490 381454
rect 266726 381218 297210 381454
rect 297446 381218 327930 381454
rect 328166 381218 358650 381454
rect 358886 381218 389370 381454
rect 389606 381218 420090 381454
rect 420326 381218 450810 381454
rect 451046 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 143610 381134
rect 143846 380898 174330 381134
rect 174566 380898 205050 381134
rect 205286 380898 235770 381134
rect 236006 380898 266490 381134
rect 266726 380898 297210 381134
rect 297446 380898 327930 381134
rect 328166 380898 358650 381134
rect 358886 380898 389370 381134
rect 389606 380898 420090 381134
rect 420326 380898 450810 381134
rect 451046 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 128250 363454
rect 128486 363218 158970 363454
rect 159206 363218 189690 363454
rect 189926 363218 220410 363454
rect 220646 363218 251130 363454
rect 251366 363218 281850 363454
rect 282086 363218 312570 363454
rect 312806 363218 343290 363454
rect 343526 363218 374010 363454
rect 374246 363218 404730 363454
rect 404966 363218 435450 363454
rect 435686 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 128250 363134
rect 128486 362898 158970 363134
rect 159206 362898 189690 363134
rect 189926 362898 220410 363134
rect 220646 362898 251130 363134
rect 251366 362898 281850 363134
rect 282086 362898 312570 363134
rect 312806 362898 343290 363134
rect 343526 362898 374010 363134
rect 374246 362898 404730 363134
rect 404966 362898 435450 363134
rect 435686 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 143610 345454
rect 143846 345218 174330 345454
rect 174566 345218 205050 345454
rect 205286 345218 235770 345454
rect 236006 345218 266490 345454
rect 266726 345218 297210 345454
rect 297446 345218 327930 345454
rect 328166 345218 358650 345454
rect 358886 345218 389370 345454
rect 389606 345218 420090 345454
rect 420326 345218 450810 345454
rect 451046 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 143610 345134
rect 143846 344898 174330 345134
rect 174566 344898 205050 345134
rect 205286 344898 235770 345134
rect 236006 344898 266490 345134
rect 266726 344898 297210 345134
rect 297446 344898 327930 345134
rect 328166 344898 358650 345134
rect 358886 344898 389370 345134
rect 389606 344898 420090 345134
rect 420326 344898 450810 345134
rect 451046 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 128250 327454
rect 128486 327218 158970 327454
rect 159206 327218 189690 327454
rect 189926 327218 220410 327454
rect 220646 327218 251130 327454
rect 251366 327218 281850 327454
rect 282086 327218 312570 327454
rect 312806 327218 343290 327454
rect 343526 327218 374010 327454
rect 374246 327218 404730 327454
rect 404966 327218 435450 327454
rect 435686 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 128250 327134
rect 128486 326898 158970 327134
rect 159206 326898 189690 327134
rect 189926 326898 220410 327134
rect 220646 326898 251130 327134
rect 251366 326898 281850 327134
rect 282086 326898 312570 327134
rect 312806 326898 343290 327134
rect 343526 326898 374010 327134
rect 374246 326898 404730 327134
rect 404966 326898 435450 327134
rect 435686 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 143610 309454
rect 143846 309218 174330 309454
rect 174566 309218 205050 309454
rect 205286 309218 235770 309454
rect 236006 309218 266490 309454
rect 266726 309218 297210 309454
rect 297446 309218 327930 309454
rect 328166 309218 358650 309454
rect 358886 309218 389370 309454
rect 389606 309218 420090 309454
rect 420326 309218 450810 309454
rect 451046 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 143610 309134
rect 143846 308898 174330 309134
rect 174566 308898 205050 309134
rect 205286 308898 235770 309134
rect 236006 308898 266490 309134
rect 266726 308898 297210 309134
rect 297446 308898 327930 309134
rect 328166 308898 358650 309134
rect 358886 308898 389370 309134
rect 389606 308898 420090 309134
rect 420326 308898 450810 309134
rect 451046 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 128250 291454
rect 128486 291218 158970 291454
rect 159206 291218 189690 291454
rect 189926 291218 220410 291454
rect 220646 291218 251130 291454
rect 251366 291218 281850 291454
rect 282086 291218 312570 291454
rect 312806 291218 343290 291454
rect 343526 291218 374010 291454
rect 374246 291218 404730 291454
rect 404966 291218 435450 291454
rect 435686 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 128250 291134
rect 128486 290898 158970 291134
rect 159206 290898 189690 291134
rect 189926 290898 220410 291134
rect 220646 290898 251130 291134
rect 251366 290898 281850 291134
rect 282086 290898 312570 291134
rect 312806 290898 343290 291134
rect 343526 290898 374010 291134
rect 374246 290898 404730 291134
rect 404966 290898 435450 291134
rect 435686 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 143610 273454
rect 143846 273218 174330 273454
rect 174566 273218 205050 273454
rect 205286 273218 235770 273454
rect 236006 273218 266490 273454
rect 266726 273218 297210 273454
rect 297446 273218 327930 273454
rect 328166 273218 358650 273454
rect 358886 273218 389370 273454
rect 389606 273218 420090 273454
rect 420326 273218 450810 273454
rect 451046 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 143610 273134
rect 143846 272898 174330 273134
rect 174566 272898 205050 273134
rect 205286 272898 235770 273134
rect 236006 272898 266490 273134
rect 266726 272898 297210 273134
rect 297446 272898 327930 273134
rect 328166 272898 358650 273134
rect 358886 272898 389370 273134
rect 389606 272898 420090 273134
rect 420326 272898 450810 273134
rect 451046 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 128250 255454
rect 128486 255218 158970 255454
rect 159206 255218 189690 255454
rect 189926 255218 220410 255454
rect 220646 255218 251130 255454
rect 251366 255218 281850 255454
rect 282086 255218 312570 255454
rect 312806 255218 343290 255454
rect 343526 255218 374010 255454
rect 374246 255218 404730 255454
rect 404966 255218 435450 255454
rect 435686 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 128250 255134
rect 128486 254898 158970 255134
rect 159206 254898 189690 255134
rect 189926 254898 220410 255134
rect 220646 254898 251130 255134
rect 251366 254898 281850 255134
rect 282086 254898 312570 255134
rect 312806 254898 343290 255134
rect 343526 254898 374010 255134
rect 374246 254898 404730 255134
rect 404966 254898 435450 255134
rect 435686 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 143610 237454
rect 143846 237218 174330 237454
rect 174566 237218 205050 237454
rect 205286 237218 235770 237454
rect 236006 237218 266490 237454
rect 266726 237218 297210 237454
rect 297446 237218 327930 237454
rect 328166 237218 358650 237454
rect 358886 237218 389370 237454
rect 389606 237218 420090 237454
rect 420326 237218 450810 237454
rect 451046 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 143610 237134
rect 143846 236898 174330 237134
rect 174566 236898 205050 237134
rect 205286 236898 235770 237134
rect 236006 236898 266490 237134
rect 266726 236898 297210 237134
rect 297446 236898 327930 237134
rect 328166 236898 358650 237134
rect 358886 236898 389370 237134
rect 389606 236898 420090 237134
rect 420326 236898 450810 237134
rect 451046 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 128250 219454
rect 128486 219218 158970 219454
rect 159206 219218 189690 219454
rect 189926 219218 220410 219454
rect 220646 219218 251130 219454
rect 251366 219218 281850 219454
rect 282086 219218 312570 219454
rect 312806 219218 343290 219454
rect 343526 219218 374010 219454
rect 374246 219218 404730 219454
rect 404966 219218 435450 219454
rect 435686 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 128250 219134
rect 128486 218898 158970 219134
rect 159206 218898 189690 219134
rect 189926 218898 220410 219134
rect 220646 218898 251130 219134
rect 251366 218898 281850 219134
rect 282086 218898 312570 219134
rect 312806 218898 343290 219134
rect 343526 218898 374010 219134
rect 374246 218898 404730 219134
rect 404966 218898 435450 219134
rect 435686 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 143610 201454
rect 143846 201218 174330 201454
rect 174566 201218 205050 201454
rect 205286 201218 235770 201454
rect 236006 201218 266490 201454
rect 266726 201218 297210 201454
rect 297446 201218 327930 201454
rect 328166 201218 358650 201454
rect 358886 201218 389370 201454
rect 389606 201218 420090 201454
rect 420326 201218 450810 201454
rect 451046 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 143610 201134
rect 143846 200898 174330 201134
rect 174566 200898 205050 201134
rect 205286 200898 235770 201134
rect 236006 200898 266490 201134
rect 266726 200898 297210 201134
rect 297446 200898 327930 201134
rect 328166 200898 358650 201134
rect 358886 200898 389370 201134
rect 389606 200898 420090 201134
rect 420326 200898 450810 201134
rect 451046 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 128250 183454
rect 128486 183218 158970 183454
rect 159206 183218 189690 183454
rect 189926 183218 220410 183454
rect 220646 183218 251130 183454
rect 251366 183218 281850 183454
rect 282086 183218 312570 183454
rect 312806 183218 343290 183454
rect 343526 183218 374010 183454
rect 374246 183218 404730 183454
rect 404966 183218 435450 183454
rect 435686 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 128250 183134
rect 128486 182898 158970 183134
rect 159206 182898 189690 183134
rect 189926 182898 220410 183134
rect 220646 182898 251130 183134
rect 251366 182898 281850 183134
rect 282086 182898 312570 183134
rect 312806 182898 343290 183134
rect 343526 182898 374010 183134
rect 374246 182898 404730 183134
rect 404966 182898 435450 183134
rect 435686 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 143610 165454
rect 143846 165218 174330 165454
rect 174566 165218 205050 165454
rect 205286 165218 235770 165454
rect 236006 165218 266490 165454
rect 266726 165218 297210 165454
rect 297446 165218 327930 165454
rect 328166 165218 358650 165454
rect 358886 165218 389370 165454
rect 389606 165218 420090 165454
rect 420326 165218 450810 165454
rect 451046 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 143610 165134
rect 143846 164898 174330 165134
rect 174566 164898 205050 165134
rect 205286 164898 235770 165134
rect 236006 164898 266490 165134
rect 266726 164898 297210 165134
rect 297446 164898 327930 165134
rect 328166 164898 358650 165134
rect 358886 164898 389370 165134
rect 389606 164898 420090 165134
rect 420326 164898 450810 165134
rect 451046 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_project  mprj
timestamp 1640967747
transform 1 0 124000 0 1 150400
box 290 0 337902 407623
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 148400 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 148400 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 148400 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 148400 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 148400 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 148400 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 148400 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 148400 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 148400 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 560023 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 560023 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 560023 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 560023 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 560023 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 560023 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 560023 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 560023 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 560023 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 148400 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 148400 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 148400 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 148400 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 148400 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 148400 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 148400 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 148400 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 148400 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 560023 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 560023 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 560023 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 560023 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 560023 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 560023 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 560023 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 560023 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 560023 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 148400 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 148400 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 148400 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 148400 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 148400 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 148400 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 148400 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 148400 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 148400 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 560023 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 560023 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 560023 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 560023 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 560023 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 560023 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 560023 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 560023 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 560023 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 148400 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 148400 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 148400 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 148400 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 148400 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 148400 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 148400 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 148400 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 148400 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 560023 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 560023 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 560023 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 560023 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 560023 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 560023 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 560023 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 560023 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 560023 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 148400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 148400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 148400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 148400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 148400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 148400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 148400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 148400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 148400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 148400 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 560023 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 560023 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 560023 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 560023 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 560023 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 560023 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 560023 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 560023 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 560023 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 560023 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 148400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 148400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 148400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 148400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 148400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 148400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 148400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 148400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 148400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 148400 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 560023 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 560023 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 560023 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 560023 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 560023 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 560023 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 560023 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 560023 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 560023 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 560023 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 148400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 148400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 148400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 148400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 148400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 148400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 148400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 148400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 148400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 148400 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 560023 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 560023 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 560023 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 560023 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 560023 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 560023 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 560023 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 560023 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 560023 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 560023 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 148400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 148400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 148400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 148400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 148400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 148400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 148400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 148400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 148400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 148400 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 560023 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 560023 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 560023 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 560023 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 560023 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 560023 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 560023 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 560023 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 560023 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 560023 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
