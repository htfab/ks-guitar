magic
tech sky130A
magscale 1 2
timestamp 1640964199
<< obsli1 >>
rect 1104 1241 337243 405297
<< obsm1 >>
rect 290 1235 337902 405680
<< metal2 >>
rect 1490 406823 1546 407623
rect 4434 406823 4490 407623
rect 7378 406823 7434 407623
rect 10322 406823 10378 407623
rect 13358 406823 13414 407623
rect 16302 406823 16358 407623
rect 19246 406823 19302 407623
rect 22190 406823 22246 407623
rect 25226 406823 25282 407623
rect 28170 406823 28226 407623
rect 31114 406823 31170 407623
rect 34058 406823 34114 407623
rect 37094 406823 37150 407623
rect 40038 406823 40094 407623
rect 42982 406823 43038 407623
rect 45926 406823 45982 407623
rect 48962 406823 49018 407623
rect 51906 406823 51962 407623
rect 54850 406823 54906 407623
rect 57794 406823 57850 407623
rect 60830 406823 60886 407623
rect 63774 406823 63830 407623
rect 66718 406823 66774 407623
rect 69662 406823 69718 407623
rect 72698 406823 72754 407623
rect 75642 406823 75698 407623
rect 78586 406823 78642 407623
rect 81530 406823 81586 407623
rect 84566 406823 84622 407623
rect 87510 406823 87566 407623
rect 90454 406823 90510 407623
rect 93398 406823 93454 407623
rect 96434 406823 96490 407623
rect 99378 406823 99434 407623
rect 102322 406823 102378 407623
rect 105266 406823 105322 407623
rect 108302 406823 108358 407623
rect 111246 406823 111302 407623
rect 114190 406823 114246 407623
rect 117134 406823 117190 407623
rect 120170 406823 120226 407623
rect 123114 406823 123170 407623
rect 126058 406823 126114 407623
rect 129002 406823 129058 407623
rect 132038 406823 132094 407623
rect 134982 406823 135038 407623
rect 137926 406823 137982 407623
rect 140870 406823 140926 407623
rect 143906 406823 143962 407623
rect 146850 406823 146906 407623
rect 149794 406823 149850 407623
rect 152738 406823 152794 407623
rect 155774 406823 155830 407623
rect 158718 406823 158774 407623
rect 161662 406823 161718 407623
rect 164606 406823 164662 407623
rect 167642 406823 167698 407623
rect 170586 406823 170642 407623
rect 173530 406823 173586 407623
rect 176566 406823 176622 407623
rect 179510 406823 179566 407623
rect 182454 406823 182510 407623
rect 185398 406823 185454 407623
rect 188434 406823 188490 407623
rect 191378 406823 191434 407623
rect 194322 406823 194378 407623
rect 197266 406823 197322 407623
rect 200302 406823 200358 407623
rect 203246 406823 203302 407623
rect 206190 406823 206246 407623
rect 209134 406823 209190 407623
rect 212170 406823 212226 407623
rect 215114 406823 215170 407623
rect 218058 406823 218114 407623
rect 221002 406823 221058 407623
rect 224038 406823 224094 407623
rect 226982 406823 227038 407623
rect 229926 406823 229982 407623
rect 232870 406823 232926 407623
rect 235906 406823 235962 407623
rect 238850 406823 238906 407623
rect 241794 406823 241850 407623
rect 244738 406823 244794 407623
rect 247774 406823 247830 407623
rect 250718 406823 250774 407623
rect 253662 406823 253718 407623
rect 256606 406823 256662 407623
rect 259642 406823 259698 407623
rect 262586 406823 262642 407623
rect 265530 406823 265586 407623
rect 268474 406823 268530 407623
rect 271510 406823 271566 407623
rect 274454 406823 274510 407623
rect 277398 406823 277454 407623
rect 280342 406823 280398 407623
rect 283378 406823 283434 407623
rect 286322 406823 286378 407623
rect 289266 406823 289322 407623
rect 292210 406823 292266 407623
rect 295246 406823 295302 407623
rect 298190 406823 298246 407623
rect 301134 406823 301190 407623
rect 304078 406823 304134 407623
rect 307114 406823 307170 407623
rect 310058 406823 310114 407623
rect 313002 406823 313058 407623
rect 315946 406823 316002 407623
rect 318982 406823 319038 407623
rect 321926 406823 321982 407623
rect 324870 406823 324926 407623
rect 327814 406823 327870 407623
rect 330850 406823 330906 407623
rect 333794 406823 333850 407623
rect 336738 406823 336794 407623
rect 294 0 350 800
rect 938 0 994 800
rect 1582 0 1638 800
rect 2318 0 2374 800
rect 2962 0 3018 800
rect 3698 0 3754 800
rect 4342 0 4398 800
rect 5078 0 5134 800
rect 5722 0 5778 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7838 0 7894 800
rect 8482 0 8538 800
rect 9126 0 9182 800
rect 9862 0 9918 800
rect 10506 0 10562 800
rect 11242 0 11298 800
rect 11886 0 11942 800
rect 12622 0 12678 800
rect 13266 0 13322 800
rect 14002 0 14058 800
rect 14646 0 14702 800
rect 15382 0 15438 800
rect 16026 0 16082 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18786 0 18842 800
rect 19430 0 19486 800
rect 20166 0 20222 800
rect 20810 0 20866 800
rect 21546 0 21602 800
rect 22190 0 22246 800
rect 22926 0 22982 800
rect 23570 0 23626 800
rect 24306 0 24362 800
rect 24950 0 25006 800
rect 25594 0 25650 800
rect 26330 0 26386 800
rect 26974 0 27030 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 29090 0 29146 800
rect 29734 0 29790 800
rect 30470 0 30526 800
rect 31114 0 31170 800
rect 31850 0 31906 800
rect 32494 0 32550 800
rect 33230 0 33286 800
rect 33874 0 33930 800
rect 34518 0 34574 800
rect 35254 0 35310 800
rect 35898 0 35954 800
rect 36634 0 36690 800
rect 37278 0 37334 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39394 0 39450 800
rect 40038 0 40094 800
rect 40774 0 40830 800
rect 41418 0 41474 800
rect 42062 0 42118 800
rect 42798 0 42854 800
rect 43442 0 43498 800
rect 44178 0 44234 800
rect 44822 0 44878 800
rect 45558 0 45614 800
rect 46202 0 46258 800
rect 46938 0 46994 800
rect 47582 0 47638 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49698 0 49754 800
rect 50342 0 50398 800
rect 50986 0 51042 800
rect 51722 0 51778 800
rect 52366 0 52422 800
rect 53102 0 53158 800
rect 53746 0 53802 800
rect 54482 0 54538 800
rect 55126 0 55182 800
rect 55862 0 55918 800
rect 56506 0 56562 800
rect 57242 0 57298 800
rect 57886 0 57942 800
rect 58530 0 58586 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 60646 0 60702 800
rect 61290 0 61346 800
rect 62026 0 62082 800
rect 62670 0 62726 800
rect 63406 0 63462 800
rect 64050 0 64106 800
rect 64786 0 64842 800
rect 65430 0 65486 800
rect 66166 0 66222 800
rect 66810 0 66866 800
rect 67454 0 67510 800
rect 68190 0 68246 800
rect 68834 0 68890 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 70950 0 71006 800
rect 71594 0 71650 800
rect 72330 0 72386 800
rect 72974 0 73030 800
rect 73710 0 73766 800
rect 74354 0 74410 800
rect 74998 0 75054 800
rect 75734 0 75790 800
rect 76378 0 76434 800
rect 77114 0 77170 800
rect 77758 0 77814 800
rect 78494 0 78550 800
rect 79138 0 79194 800
rect 79874 0 79930 800
rect 80518 0 80574 800
rect 81254 0 81310 800
rect 81898 0 81954 800
rect 82634 0 82690 800
rect 83278 0 83334 800
rect 83922 0 83978 800
rect 84658 0 84714 800
rect 85302 0 85358 800
rect 86038 0 86094 800
rect 86682 0 86738 800
rect 87418 0 87474 800
rect 88062 0 88118 800
rect 88798 0 88854 800
rect 89442 0 89498 800
rect 90178 0 90234 800
rect 90822 0 90878 800
rect 91466 0 91522 800
rect 92202 0 92258 800
rect 92846 0 92902 800
rect 93582 0 93638 800
rect 94226 0 94282 800
rect 94962 0 95018 800
rect 95606 0 95662 800
rect 96342 0 96398 800
rect 96986 0 97042 800
rect 97722 0 97778 800
rect 98366 0 98422 800
rect 99102 0 99158 800
rect 99746 0 99802 800
rect 100390 0 100446 800
rect 101126 0 101182 800
rect 101770 0 101826 800
rect 102506 0 102562 800
rect 103150 0 103206 800
rect 103886 0 103942 800
rect 104530 0 104586 800
rect 105266 0 105322 800
rect 105910 0 105966 800
rect 106646 0 106702 800
rect 107290 0 107346 800
rect 107934 0 107990 800
rect 108670 0 108726 800
rect 109314 0 109370 800
rect 110050 0 110106 800
rect 110694 0 110750 800
rect 111430 0 111486 800
rect 112074 0 112130 800
rect 112810 0 112866 800
rect 113454 0 113510 800
rect 114190 0 114246 800
rect 114834 0 114890 800
rect 115570 0 115626 800
rect 116214 0 116270 800
rect 116858 0 116914 800
rect 117594 0 117650 800
rect 118238 0 118294 800
rect 118974 0 119030 800
rect 119618 0 119674 800
rect 120354 0 120410 800
rect 120998 0 121054 800
rect 121734 0 121790 800
rect 122378 0 122434 800
rect 123114 0 123170 800
rect 123758 0 123814 800
rect 124402 0 124458 800
rect 125138 0 125194 800
rect 125782 0 125838 800
rect 126518 0 126574 800
rect 127162 0 127218 800
rect 127898 0 127954 800
rect 128542 0 128598 800
rect 129278 0 129334 800
rect 129922 0 129978 800
rect 130658 0 130714 800
rect 131302 0 131358 800
rect 132038 0 132094 800
rect 132682 0 132738 800
rect 133326 0 133382 800
rect 134062 0 134118 800
rect 134706 0 134762 800
rect 135442 0 135498 800
rect 136086 0 136142 800
rect 136822 0 136878 800
rect 137466 0 137522 800
rect 138202 0 138258 800
rect 138846 0 138902 800
rect 139582 0 139638 800
rect 140226 0 140282 800
rect 140870 0 140926 800
rect 141606 0 141662 800
rect 142250 0 142306 800
rect 142986 0 143042 800
rect 143630 0 143686 800
rect 144366 0 144422 800
rect 145010 0 145066 800
rect 145746 0 145802 800
rect 146390 0 146446 800
rect 147126 0 147182 800
rect 147770 0 147826 800
rect 148506 0 148562 800
rect 149150 0 149206 800
rect 149794 0 149850 800
rect 150530 0 150586 800
rect 151174 0 151230 800
rect 151910 0 151966 800
rect 152554 0 152610 800
rect 153290 0 153346 800
rect 153934 0 153990 800
rect 154670 0 154726 800
rect 155314 0 155370 800
rect 156050 0 156106 800
rect 156694 0 156750 800
rect 157338 0 157394 800
rect 158074 0 158130 800
rect 158718 0 158774 800
rect 159454 0 159510 800
rect 160098 0 160154 800
rect 160834 0 160890 800
rect 161478 0 161534 800
rect 162214 0 162270 800
rect 162858 0 162914 800
rect 163594 0 163650 800
rect 164238 0 164294 800
rect 164974 0 165030 800
rect 165618 0 165674 800
rect 166262 0 166318 800
rect 166998 0 167054 800
rect 167642 0 167698 800
rect 168378 0 168434 800
rect 169022 0 169078 800
rect 169758 0 169814 800
rect 170402 0 170458 800
rect 171138 0 171194 800
rect 171782 0 171838 800
rect 172518 0 172574 800
rect 173162 0 173218 800
rect 173806 0 173862 800
rect 174542 0 174598 800
rect 175186 0 175242 800
rect 175922 0 175978 800
rect 176566 0 176622 800
rect 177302 0 177358 800
rect 177946 0 178002 800
rect 178682 0 178738 800
rect 179326 0 179382 800
rect 180062 0 180118 800
rect 180706 0 180762 800
rect 181442 0 181498 800
rect 182086 0 182142 800
rect 182730 0 182786 800
rect 183466 0 183522 800
rect 184110 0 184166 800
rect 184846 0 184902 800
rect 185490 0 185546 800
rect 186226 0 186282 800
rect 186870 0 186926 800
rect 187606 0 187662 800
rect 188250 0 188306 800
rect 188986 0 189042 800
rect 189630 0 189686 800
rect 190274 0 190330 800
rect 191010 0 191066 800
rect 191654 0 191710 800
rect 192390 0 192446 800
rect 193034 0 193090 800
rect 193770 0 193826 800
rect 194414 0 194470 800
rect 195150 0 195206 800
rect 195794 0 195850 800
rect 196530 0 196586 800
rect 197174 0 197230 800
rect 197910 0 197966 800
rect 198554 0 198610 800
rect 199198 0 199254 800
rect 199934 0 199990 800
rect 200578 0 200634 800
rect 201314 0 201370 800
rect 201958 0 202014 800
rect 202694 0 202750 800
rect 203338 0 203394 800
rect 204074 0 204130 800
rect 204718 0 204774 800
rect 205454 0 205510 800
rect 206098 0 206154 800
rect 206742 0 206798 800
rect 207478 0 207534 800
rect 208122 0 208178 800
rect 208858 0 208914 800
rect 209502 0 209558 800
rect 210238 0 210294 800
rect 210882 0 210938 800
rect 211618 0 211674 800
rect 212262 0 212318 800
rect 212998 0 213054 800
rect 213642 0 213698 800
rect 214378 0 214434 800
rect 215022 0 215078 800
rect 215666 0 215722 800
rect 216402 0 216458 800
rect 217046 0 217102 800
rect 217782 0 217838 800
rect 218426 0 218482 800
rect 219162 0 219218 800
rect 219806 0 219862 800
rect 220542 0 220598 800
rect 221186 0 221242 800
rect 221922 0 221978 800
rect 222566 0 222622 800
rect 223210 0 223266 800
rect 223946 0 224002 800
rect 224590 0 224646 800
rect 225326 0 225382 800
rect 225970 0 226026 800
rect 226706 0 226762 800
rect 227350 0 227406 800
rect 228086 0 228142 800
rect 228730 0 228786 800
rect 229466 0 229522 800
rect 230110 0 230166 800
rect 230846 0 230902 800
rect 231490 0 231546 800
rect 232134 0 232190 800
rect 232870 0 232926 800
rect 233514 0 233570 800
rect 234250 0 234306 800
rect 234894 0 234950 800
rect 235630 0 235686 800
rect 236274 0 236330 800
rect 237010 0 237066 800
rect 237654 0 237710 800
rect 238390 0 238446 800
rect 239034 0 239090 800
rect 239678 0 239734 800
rect 240414 0 240470 800
rect 241058 0 241114 800
rect 241794 0 241850 800
rect 242438 0 242494 800
rect 243174 0 243230 800
rect 243818 0 243874 800
rect 244554 0 244610 800
rect 245198 0 245254 800
rect 245934 0 245990 800
rect 246578 0 246634 800
rect 247314 0 247370 800
rect 247958 0 248014 800
rect 248602 0 248658 800
rect 249338 0 249394 800
rect 249982 0 250038 800
rect 250718 0 250774 800
rect 251362 0 251418 800
rect 252098 0 252154 800
rect 252742 0 252798 800
rect 253478 0 253534 800
rect 254122 0 254178 800
rect 254858 0 254914 800
rect 255502 0 255558 800
rect 256146 0 256202 800
rect 256882 0 256938 800
rect 257526 0 257582 800
rect 258262 0 258318 800
rect 258906 0 258962 800
rect 259642 0 259698 800
rect 260286 0 260342 800
rect 261022 0 261078 800
rect 261666 0 261722 800
rect 262402 0 262458 800
rect 263046 0 263102 800
rect 263782 0 263838 800
rect 264426 0 264482 800
rect 265070 0 265126 800
rect 265806 0 265862 800
rect 266450 0 266506 800
rect 267186 0 267242 800
rect 267830 0 267886 800
rect 268566 0 268622 800
rect 269210 0 269266 800
rect 269946 0 270002 800
rect 270590 0 270646 800
rect 271326 0 271382 800
rect 271970 0 272026 800
rect 272614 0 272670 800
rect 273350 0 273406 800
rect 273994 0 274050 800
rect 274730 0 274786 800
rect 275374 0 275430 800
rect 276110 0 276166 800
rect 276754 0 276810 800
rect 277490 0 277546 800
rect 278134 0 278190 800
rect 278870 0 278926 800
rect 279514 0 279570 800
rect 280250 0 280306 800
rect 280894 0 280950 800
rect 281538 0 281594 800
rect 282274 0 282330 800
rect 282918 0 282974 800
rect 283654 0 283710 800
rect 284298 0 284354 800
rect 285034 0 285090 800
rect 285678 0 285734 800
rect 286414 0 286470 800
rect 287058 0 287114 800
rect 287794 0 287850 800
rect 288438 0 288494 800
rect 289082 0 289138 800
rect 289818 0 289874 800
rect 290462 0 290518 800
rect 291198 0 291254 800
rect 291842 0 291898 800
rect 292578 0 292634 800
rect 293222 0 293278 800
rect 293958 0 294014 800
rect 294602 0 294658 800
rect 295338 0 295394 800
rect 295982 0 296038 800
rect 296718 0 296774 800
rect 297362 0 297418 800
rect 298006 0 298062 800
rect 298742 0 298798 800
rect 299386 0 299442 800
rect 300122 0 300178 800
rect 300766 0 300822 800
rect 301502 0 301558 800
rect 302146 0 302202 800
rect 302882 0 302938 800
rect 303526 0 303582 800
rect 304262 0 304318 800
rect 304906 0 304962 800
rect 305550 0 305606 800
rect 306286 0 306342 800
rect 306930 0 306986 800
rect 307666 0 307722 800
rect 308310 0 308366 800
rect 309046 0 309102 800
rect 309690 0 309746 800
rect 310426 0 310482 800
rect 311070 0 311126 800
rect 311806 0 311862 800
rect 312450 0 312506 800
rect 313186 0 313242 800
rect 313830 0 313886 800
rect 314474 0 314530 800
rect 315210 0 315266 800
rect 315854 0 315910 800
rect 316590 0 316646 800
rect 317234 0 317290 800
rect 317970 0 318026 800
rect 318614 0 318670 800
rect 319350 0 319406 800
rect 319994 0 320050 800
rect 320730 0 320786 800
rect 321374 0 321430 800
rect 322018 0 322074 800
rect 322754 0 322810 800
rect 323398 0 323454 800
rect 324134 0 324190 800
rect 324778 0 324834 800
rect 325514 0 325570 800
rect 326158 0 326214 800
rect 326894 0 326950 800
rect 327538 0 327594 800
rect 328274 0 328330 800
rect 328918 0 328974 800
rect 329654 0 329710 800
rect 330298 0 330354 800
rect 330942 0 330998 800
rect 331678 0 331734 800
rect 332322 0 332378 800
rect 333058 0 333114 800
rect 333702 0 333758 800
rect 334438 0 334494 800
rect 335082 0 335138 800
rect 335818 0 335874 800
rect 336462 0 336518 800
rect 337198 0 337254 800
rect 337842 0 337898 800
<< obsm2 >>
rect 296 406767 1434 406858
rect 1602 406767 4378 406858
rect 4546 406767 7322 406858
rect 7490 406767 10266 406858
rect 10434 406767 13302 406858
rect 13470 406767 16246 406858
rect 16414 406767 19190 406858
rect 19358 406767 22134 406858
rect 22302 406767 25170 406858
rect 25338 406767 28114 406858
rect 28282 406767 31058 406858
rect 31226 406767 34002 406858
rect 34170 406767 37038 406858
rect 37206 406767 39982 406858
rect 40150 406767 42926 406858
rect 43094 406767 45870 406858
rect 46038 406767 48906 406858
rect 49074 406767 51850 406858
rect 52018 406767 54794 406858
rect 54962 406767 57738 406858
rect 57906 406767 60774 406858
rect 60942 406767 63718 406858
rect 63886 406767 66662 406858
rect 66830 406767 69606 406858
rect 69774 406767 72642 406858
rect 72810 406767 75586 406858
rect 75754 406767 78530 406858
rect 78698 406767 81474 406858
rect 81642 406767 84510 406858
rect 84678 406767 87454 406858
rect 87622 406767 90398 406858
rect 90566 406767 93342 406858
rect 93510 406767 96378 406858
rect 96546 406767 99322 406858
rect 99490 406767 102266 406858
rect 102434 406767 105210 406858
rect 105378 406767 108246 406858
rect 108414 406767 111190 406858
rect 111358 406767 114134 406858
rect 114302 406767 117078 406858
rect 117246 406767 120114 406858
rect 120282 406767 123058 406858
rect 123226 406767 126002 406858
rect 126170 406767 128946 406858
rect 129114 406767 131982 406858
rect 132150 406767 134926 406858
rect 135094 406767 137870 406858
rect 138038 406767 140814 406858
rect 140982 406767 143850 406858
rect 144018 406767 146794 406858
rect 146962 406767 149738 406858
rect 149906 406767 152682 406858
rect 152850 406767 155718 406858
rect 155886 406767 158662 406858
rect 158830 406767 161606 406858
rect 161774 406767 164550 406858
rect 164718 406767 167586 406858
rect 167754 406767 170530 406858
rect 170698 406767 173474 406858
rect 173642 406767 176510 406858
rect 176678 406767 179454 406858
rect 179622 406767 182398 406858
rect 182566 406767 185342 406858
rect 185510 406767 188378 406858
rect 188546 406767 191322 406858
rect 191490 406767 194266 406858
rect 194434 406767 197210 406858
rect 197378 406767 200246 406858
rect 200414 406767 203190 406858
rect 203358 406767 206134 406858
rect 206302 406767 209078 406858
rect 209246 406767 212114 406858
rect 212282 406767 215058 406858
rect 215226 406767 218002 406858
rect 218170 406767 220946 406858
rect 221114 406767 223982 406858
rect 224150 406767 226926 406858
rect 227094 406767 229870 406858
rect 230038 406767 232814 406858
rect 232982 406767 235850 406858
rect 236018 406767 238794 406858
rect 238962 406767 241738 406858
rect 241906 406767 244682 406858
rect 244850 406767 247718 406858
rect 247886 406767 250662 406858
rect 250830 406767 253606 406858
rect 253774 406767 256550 406858
rect 256718 406767 259586 406858
rect 259754 406767 262530 406858
rect 262698 406767 265474 406858
rect 265642 406767 268418 406858
rect 268586 406767 271454 406858
rect 271622 406767 274398 406858
rect 274566 406767 277342 406858
rect 277510 406767 280286 406858
rect 280454 406767 283322 406858
rect 283490 406767 286266 406858
rect 286434 406767 289210 406858
rect 289378 406767 292154 406858
rect 292322 406767 295190 406858
rect 295358 406767 298134 406858
rect 298302 406767 301078 406858
rect 301246 406767 304022 406858
rect 304190 406767 307058 406858
rect 307226 406767 310002 406858
rect 310170 406767 312946 406858
rect 313114 406767 315890 406858
rect 316058 406767 318926 406858
rect 319094 406767 321870 406858
rect 322038 406767 324814 406858
rect 324982 406767 327758 406858
rect 327926 406767 330794 406858
rect 330962 406767 333738 406858
rect 333906 406767 336682 406858
rect 336850 406767 337896 406858
rect 296 856 337896 406767
rect 406 734 882 856
rect 1050 734 1526 856
rect 1694 734 2262 856
rect 2430 734 2906 856
rect 3074 734 3642 856
rect 3810 734 4286 856
rect 4454 734 5022 856
rect 5190 734 5666 856
rect 5834 734 6402 856
rect 6570 734 7046 856
rect 7214 734 7782 856
rect 7950 734 8426 856
rect 8594 734 9070 856
rect 9238 734 9806 856
rect 9974 734 10450 856
rect 10618 734 11186 856
rect 11354 734 11830 856
rect 11998 734 12566 856
rect 12734 734 13210 856
rect 13378 734 13946 856
rect 14114 734 14590 856
rect 14758 734 15326 856
rect 15494 734 15970 856
rect 16138 734 16706 856
rect 16874 734 17350 856
rect 17518 734 17994 856
rect 18162 734 18730 856
rect 18898 734 19374 856
rect 19542 734 20110 856
rect 20278 734 20754 856
rect 20922 734 21490 856
rect 21658 734 22134 856
rect 22302 734 22870 856
rect 23038 734 23514 856
rect 23682 734 24250 856
rect 24418 734 24894 856
rect 25062 734 25538 856
rect 25706 734 26274 856
rect 26442 734 26918 856
rect 27086 734 27654 856
rect 27822 734 28298 856
rect 28466 734 29034 856
rect 29202 734 29678 856
rect 29846 734 30414 856
rect 30582 734 31058 856
rect 31226 734 31794 856
rect 31962 734 32438 856
rect 32606 734 33174 856
rect 33342 734 33818 856
rect 33986 734 34462 856
rect 34630 734 35198 856
rect 35366 734 35842 856
rect 36010 734 36578 856
rect 36746 734 37222 856
rect 37390 734 37958 856
rect 38126 734 38602 856
rect 38770 734 39338 856
rect 39506 734 39982 856
rect 40150 734 40718 856
rect 40886 734 41362 856
rect 41530 734 42006 856
rect 42174 734 42742 856
rect 42910 734 43386 856
rect 43554 734 44122 856
rect 44290 734 44766 856
rect 44934 734 45502 856
rect 45670 734 46146 856
rect 46314 734 46882 856
rect 47050 734 47526 856
rect 47694 734 48262 856
rect 48430 734 48906 856
rect 49074 734 49642 856
rect 49810 734 50286 856
rect 50454 734 50930 856
rect 51098 734 51666 856
rect 51834 734 52310 856
rect 52478 734 53046 856
rect 53214 734 53690 856
rect 53858 734 54426 856
rect 54594 734 55070 856
rect 55238 734 55806 856
rect 55974 734 56450 856
rect 56618 734 57186 856
rect 57354 734 57830 856
rect 57998 734 58474 856
rect 58642 734 59210 856
rect 59378 734 59854 856
rect 60022 734 60590 856
rect 60758 734 61234 856
rect 61402 734 61970 856
rect 62138 734 62614 856
rect 62782 734 63350 856
rect 63518 734 63994 856
rect 64162 734 64730 856
rect 64898 734 65374 856
rect 65542 734 66110 856
rect 66278 734 66754 856
rect 66922 734 67398 856
rect 67566 734 68134 856
rect 68302 734 68778 856
rect 68946 734 69514 856
rect 69682 734 70158 856
rect 70326 734 70894 856
rect 71062 734 71538 856
rect 71706 734 72274 856
rect 72442 734 72918 856
rect 73086 734 73654 856
rect 73822 734 74298 856
rect 74466 734 74942 856
rect 75110 734 75678 856
rect 75846 734 76322 856
rect 76490 734 77058 856
rect 77226 734 77702 856
rect 77870 734 78438 856
rect 78606 734 79082 856
rect 79250 734 79818 856
rect 79986 734 80462 856
rect 80630 734 81198 856
rect 81366 734 81842 856
rect 82010 734 82578 856
rect 82746 734 83222 856
rect 83390 734 83866 856
rect 84034 734 84602 856
rect 84770 734 85246 856
rect 85414 734 85982 856
rect 86150 734 86626 856
rect 86794 734 87362 856
rect 87530 734 88006 856
rect 88174 734 88742 856
rect 88910 734 89386 856
rect 89554 734 90122 856
rect 90290 734 90766 856
rect 90934 734 91410 856
rect 91578 734 92146 856
rect 92314 734 92790 856
rect 92958 734 93526 856
rect 93694 734 94170 856
rect 94338 734 94906 856
rect 95074 734 95550 856
rect 95718 734 96286 856
rect 96454 734 96930 856
rect 97098 734 97666 856
rect 97834 734 98310 856
rect 98478 734 99046 856
rect 99214 734 99690 856
rect 99858 734 100334 856
rect 100502 734 101070 856
rect 101238 734 101714 856
rect 101882 734 102450 856
rect 102618 734 103094 856
rect 103262 734 103830 856
rect 103998 734 104474 856
rect 104642 734 105210 856
rect 105378 734 105854 856
rect 106022 734 106590 856
rect 106758 734 107234 856
rect 107402 734 107878 856
rect 108046 734 108614 856
rect 108782 734 109258 856
rect 109426 734 109994 856
rect 110162 734 110638 856
rect 110806 734 111374 856
rect 111542 734 112018 856
rect 112186 734 112754 856
rect 112922 734 113398 856
rect 113566 734 114134 856
rect 114302 734 114778 856
rect 114946 734 115514 856
rect 115682 734 116158 856
rect 116326 734 116802 856
rect 116970 734 117538 856
rect 117706 734 118182 856
rect 118350 734 118918 856
rect 119086 734 119562 856
rect 119730 734 120298 856
rect 120466 734 120942 856
rect 121110 734 121678 856
rect 121846 734 122322 856
rect 122490 734 123058 856
rect 123226 734 123702 856
rect 123870 734 124346 856
rect 124514 734 125082 856
rect 125250 734 125726 856
rect 125894 734 126462 856
rect 126630 734 127106 856
rect 127274 734 127842 856
rect 128010 734 128486 856
rect 128654 734 129222 856
rect 129390 734 129866 856
rect 130034 734 130602 856
rect 130770 734 131246 856
rect 131414 734 131982 856
rect 132150 734 132626 856
rect 132794 734 133270 856
rect 133438 734 134006 856
rect 134174 734 134650 856
rect 134818 734 135386 856
rect 135554 734 136030 856
rect 136198 734 136766 856
rect 136934 734 137410 856
rect 137578 734 138146 856
rect 138314 734 138790 856
rect 138958 734 139526 856
rect 139694 734 140170 856
rect 140338 734 140814 856
rect 140982 734 141550 856
rect 141718 734 142194 856
rect 142362 734 142930 856
rect 143098 734 143574 856
rect 143742 734 144310 856
rect 144478 734 144954 856
rect 145122 734 145690 856
rect 145858 734 146334 856
rect 146502 734 147070 856
rect 147238 734 147714 856
rect 147882 734 148450 856
rect 148618 734 149094 856
rect 149262 734 149738 856
rect 149906 734 150474 856
rect 150642 734 151118 856
rect 151286 734 151854 856
rect 152022 734 152498 856
rect 152666 734 153234 856
rect 153402 734 153878 856
rect 154046 734 154614 856
rect 154782 734 155258 856
rect 155426 734 155994 856
rect 156162 734 156638 856
rect 156806 734 157282 856
rect 157450 734 158018 856
rect 158186 734 158662 856
rect 158830 734 159398 856
rect 159566 734 160042 856
rect 160210 734 160778 856
rect 160946 734 161422 856
rect 161590 734 162158 856
rect 162326 734 162802 856
rect 162970 734 163538 856
rect 163706 734 164182 856
rect 164350 734 164918 856
rect 165086 734 165562 856
rect 165730 734 166206 856
rect 166374 734 166942 856
rect 167110 734 167586 856
rect 167754 734 168322 856
rect 168490 734 168966 856
rect 169134 734 169702 856
rect 169870 734 170346 856
rect 170514 734 171082 856
rect 171250 734 171726 856
rect 171894 734 172462 856
rect 172630 734 173106 856
rect 173274 734 173750 856
rect 173918 734 174486 856
rect 174654 734 175130 856
rect 175298 734 175866 856
rect 176034 734 176510 856
rect 176678 734 177246 856
rect 177414 734 177890 856
rect 178058 734 178626 856
rect 178794 734 179270 856
rect 179438 734 180006 856
rect 180174 734 180650 856
rect 180818 734 181386 856
rect 181554 734 182030 856
rect 182198 734 182674 856
rect 182842 734 183410 856
rect 183578 734 184054 856
rect 184222 734 184790 856
rect 184958 734 185434 856
rect 185602 734 186170 856
rect 186338 734 186814 856
rect 186982 734 187550 856
rect 187718 734 188194 856
rect 188362 734 188930 856
rect 189098 734 189574 856
rect 189742 734 190218 856
rect 190386 734 190954 856
rect 191122 734 191598 856
rect 191766 734 192334 856
rect 192502 734 192978 856
rect 193146 734 193714 856
rect 193882 734 194358 856
rect 194526 734 195094 856
rect 195262 734 195738 856
rect 195906 734 196474 856
rect 196642 734 197118 856
rect 197286 734 197854 856
rect 198022 734 198498 856
rect 198666 734 199142 856
rect 199310 734 199878 856
rect 200046 734 200522 856
rect 200690 734 201258 856
rect 201426 734 201902 856
rect 202070 734 202638 856
rect 202806 734 203282 856
rect 203450 734 204018 856
rect 204186 734 204662 856
rect 204830 734 205398 856
rect 205566 734 206042 856
rect 206210 734 206686 856
rect 206854 734 207422 856
rect 207590 734 208066 856
rect 208234 734 208802 856
rect 208970 734 209446 856
rect 209614 734 210182 856
rect 210350 734 210826 856
rect 210994 734 211562 856
rect 211730 734 212206 856
rect 212374 734 212942 856
rect 213110 734 213586 856
rect 213754 734 214322 856
rect 214490 734 214966 856
rect 215134 734 215610 856
rect 215778 734 216346 856
rect 216514 734 216990 856
rect 217158 734 217726 856
rect 217894 734 218370 856
rect 218538 734 219106 856
rect 219274 734 219750 856
rect 219918 734 220486 856
rect 220654 734 221130 856
rect 221298 734 221866 856
rect 222034 734 222510 856
rect 222678 734 223154 856
rect 223322 734 223890 856
rect 224058 734 224534 856
rect 224702 734 225270 856
rect 225438 734 225914 856
rect 226082 734 226650 856
rect 226818 734 227294 856
rect 227462 734 228030 856
rect 228198 734 228674 856
rect 228842 734 229410 856
rect 229578 734 230054 856
rect 230222 734 230790 856
rect 230958 734 231434 856
rect 231602 734 232078 856
rect 232246 734 232814 856
rect 232982 734 233458 856
rect 233626 734 234194 856
rect 234362 734 234838 856
rect 235006 734 235574 856
rect 235742 734 236218 856
rect 236386 734 236954 856
rect 237122 734 237598 856
rect 237766 734 238334 856
rect 238502 734 238978 856
rect 239146 734 239622 856
rect 239790 734 240358 856
rect 240526 734 241002 856
rect 241170 734 241738 856
rect 241906 734 242382 856
rect 242550 734 243118 856
rect 243286 734 243762 856
rect 243930 734 244498 856
rect 244666 734 245142 856
rect 245310 734 245878 856
rect 246046 734 246522 856
rect 246690 734 247258 856
rect 247426 734 247902 856
rect 248070 734 248546 856
rect 248714 734 249282 856
rect 249450 734 249926 856
rect 250094 734 250662 856
rect 250830 734 251306 856
rect 251474 734 252042 856
rect 252210 734 252686 856
rect 252854 734 253422 856
rect 253590 734 254066 856
rect 254234 734 254802 856
rect 254970 734 255446 856
rect 255614 734 256090 856
rect 256258 734 256826 856
rect 256994 734 257470 856
rect 257638 734 258206 856
rect 258374 734 258850 856
rect 259018 734 259586 856
rect 259754 734 260230 856
rect 260398 734 260966 856
rect 261134 734 261610 856
rect 261778 734 262346 856
rect 262514 734 262990 856
rect 263158 734 263726 856
rect 263894 734 264370 856
rect 264538 734 265014 856
rect 265182 734 265750 856
rect 265918 734 266394 856
rect 266562 734 267130 856
rect 267298 734 267774 856
rect 267942 734 268510 856
rect 268678 734 269154 856
rect 269322 734 269890 856
rect 270058 734 270534 856
rect 270702 734 271270 856
rect 271438 734 271914 856
rect 272082 734 272558 856
rect 272726 734 273294 856
rect 273462 734 273938 856
rect 274106 734 274674 856
rect 274842 734 275318 856
rect 275486 734 276054 856
rect 276222 734 276698 856
rect 276866 734 277434 856
rect 277602 734 278078 856
rect 278246 734 278814 856
rect 278982 734 279458 856
rect 279626 734 280194 856
rect 280362 734 280838 856
rect 281006 734 281482 856
rect 281650 734 282218 856
rect 282386 734 282862 856
rect 283030 734 283598 856
rect 283766 734 284242 856
rect 284410 734 284978 856
rect 285146 734 285622 856
rect 285790 734 286358 856
rect 286526 734 287002 856
rect 287170 734 287738 856
rect 287906 734 288382 856
rect 288550 734 289026 856
rect 289194 734 289762 856
rect 289930 734 290406 856
rect 290574 734 291142 856
rect 291310 734 291786 856
rect 291954 734 292522 856
rect 292690 734 293166 856
rect 293334 734 293902 856
rect 294070 734 294546 856
rect 294714 734 295282 856
rect 295450 734 295926 856
rect 296094 734 296662 856
rect 296830 734 297306 856
rect 297474 734 297950 856
rect 298118 734 298686 856
rect 298854 734 299330 856
rect 299498 734 300066 856
rect 300234 734 300710 856
rect 300878 734 301446 856
rect 301614 734 302090 856
rect 302258 734 302826 856
rect 302994 734 303470 856
rect 303638 734 304206 856
rect 304374 734 304850 856
rect 305018 734 305494 856
rect 305662 734 306230 856
rect 306398 734 306874 856
rect 307042 734 307610 856
rect 307778 734 308254 856
rect 308422 734 308990 856
rect 309158 734 309634 856
rect 309802 734 310370 856
rect 310538 734 311014 856
rect 311182 734 311750 856
rect 311918 734 312394 856
rect 312562 734 313130 856
rect 313298 734 313774 856
rect 313942 734 314418 856
rect 314586 734 315154 856
rect 315322 734 315798 856
rect 315966 734 316534 856
rect 316702 734 317178 856
rect 317346 734 317914 856
rect 318082 734 318558 856
rect 318726 734 319294 856
rect 319462 734 319938 856
rect 320106 734 320674 856
rect 320842 734 321318 856
rect 321486 734 321962 856
rect 322130 734 322698 856
rect 322866 734 323342 856
rect 323510 734 324078 856
rect 324246 734 324722 856
rect 324890 734 325458 856
rect 325626 734 326102 856
rect 326270 734 326838 856
rect 327006 734 327482 856
rect 327650 734 328218 856
rect 328386 734 328862 856
rect 329030 734 329598 856
rect 329766 734 330242 856
rect 330410 734 330886 856
rect 331054 734 331622 856
rect 331790 734 332266 856
rect 332434 734 333002 856
rect 333170 734 333646 856
rect 333814 734 334382 856
rect 334550 734 335026 856
rect 335194 734 335762 856
rect 335930 734 336406 856
rect 336574 734 337142 856
rect 337310 734 337786 856
<< obsm3 >>
rect 4208 1803 331279 405313
<< metal4 >>
rect 4208 2128 4528 405328
rect 19568 2128 19888 405328
rect 34928 2128 35248 405328
rect 50288 2128 50608 405328
rect 65648 2128 65968 405328
rect 81008 2128 81328 405328
rect 96368 2128 96688 405328
rect 111728 2128 112048 405328
rect 127088 2128 127408 405328
rect 142448 2128 142768 405328
rect 157808 2128 158128 405328
rect 173168 2128 173488 405328
rect 188528 2128 188848 405328
rect 203888 2128 204208 405328
rect 219248 2128 219568 405328
rect 234608 2128 234928 405328
rect 249968 2128 250288 405328
rect 265328 2128 265648 405328
rect 280688 2128 281008 405328
rect 296048 2128 296368 405328
rect 311408 2128 311728 405328
rect 326768 2128 327088 405328
<< obsm4 >>
rect 38699 3707 50208 401709
rect 50688 3707 65568 401709
rect 66048 3707 80928 401709
rect 81408 3707 96288 401709
rect 96768 3707 111648 401709
rect 112128 3707 127008 401709
rect 127488 3707 142368 401709
rect 142848 3707 157728 401709
rect 158208 3707 173088 401709
rect 173568 3707 188448 401709
rect 188928 3707 203808 401709
rect 204288 3707 219168 401709
rect 219648 3707 234528 401709
rect 235008 3707 249888 401709
rect 250368 3707 265248 401709
rect 265728 3707 280608 401709
rect 281088 3707 295968 401709
rect 296448 3707 311269 401709
<< labels >>
rlabel metal2 s 1490 406823 1546 407623 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 90454 406823 90510 407623 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 99378 406823 99434 407623 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 108302 406823 108358 407623 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 117134 406823 117190 407623 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 126058 406823 126114 407623 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 134982 406823 135038 407623 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 143906 406823 143962 407623 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 152738 406823 152794 407623 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 161662 406823 161718 407623 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 170586 406823 170642 407623 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 10322 406823 10378 407623 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 179510 406823 179566 407623 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 188434 406823 188490 407623 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 197266 406823 197322 407623 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 206190 406823 206246 407623 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 215114 406823 215170 407623 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 224038 406823 224094 407623 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 232870 406823 232926 407623 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 241794 406823 241850 407623 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 250718 406823 250774 407623 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 259642 406823 259698 407623 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 19246 406823 19302 407623 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 268474 406823 268530 407623 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 277398 406823 277454 407623 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 286322 406823 286378 407623 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 295246 406823 295302 407623 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 304078 406823 304134 407623 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 313002 406823 313058 407623 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 321926 406823 321982 407623 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 330850 406823 330906 407623 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 28170 406823 28226 407623 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 37094 406823 37150 407623 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 45926 406823 45982 407623 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 54850 406823 54906 407623 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 63774 406823 63830 407623 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 72698 406823 72754 407623 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 81530 406823 81586 407623 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 4434 406823 4490 407623 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 93398 406823 93454 407623 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 102322 406823 102378 407623 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 111246 406823 111302 407623 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 120170 406823 120226 407623 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 129002 406823 129058 407623 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 137926 406823 137982 407623 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 146850 406823 146906 407623 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 155774 406823 155830 407623 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 164606 406823 164662 407623 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 173530 406823 173586 407623 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 13358 406823 13414 407623 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 182454 406823 182510 407623 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 191378 406823 191434 407623 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 200302 406823 200358 407623 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 209134 406823 209190 407623 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 218058 406823 218114 407623 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 226982 406823 227038 407623 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 235906 406823 235962 407623 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 244738 406823 244794 407623 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 253662 406823 253718 407623 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 262586 406823 262642 407623 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 22190 406823 22246 407623 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 271510 406823 271566 407623 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 280342 406823 280398 407623 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 289266 406823 289322 407623 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 298190 406823 298246 407623 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 307114 406823 307170 407623 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 315946 406823 316002 407623 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 324870 406823 324926 407623 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 333794 406823 333850 407623 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 31114 406823 31170 407623 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 40038 406823 40094 407623 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 48962 406823 49018 407623 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 57794 406823 57850 407623 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 66718 406823 66774 407623 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 75642 406823 75698 407623 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 84566 406823 84622 407623 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 7378 406823 7434 407623 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 96434 406823 96490 407623 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 105266 406823 105322 407623 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 114190 406823 114246 407623 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 123114 406823 123170 407623 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 132038 406823 132094 407623 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 140870 406823 140926 407623 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 149794 406823 149850 407623 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 158718 406823 158774 407623 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 167642 406823 167698 407623 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 176566 406823 176622 407623 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 16302 406823 16358 407623 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 185398 406823 185454 407623 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 194322 406823 194378 407623 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 203246 406823 203302 407623 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 212170 406823 212226 407623 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 221002 406823 221058 407623 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 229926 406823 229982 407623 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 238850 406823 238906 407623 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 247774 406823 247830 407623 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 256606 406823 256662 407623 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 265530 406823 265586 407623 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 25226 406823 25282 407623 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 274454 406823 274510 407623 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 283378 406823 283434 407623 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 292210 406823 292266 407623 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 301134 406823 301190 407623 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 310058 406823 310114 407623 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 318982 406823 319038 407623 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 327814 406823 327870 407623 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 336738 406823 336794 407623 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 34058 406823 34114 407623 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 42982 406823 43038 407623 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 51906 406823 51962 407623 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 60830 406823 60886 407623 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 69662 406823 69718 407623 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 78586 406823 78642 407623 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 87510 406823 87566 407623 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 336462 0 336518 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 337198 0 337254 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 337842 0 337898 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 72974 0 73030 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 278870 0 278926 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 280894 0 280950 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 282918 0 282974 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 285034 0 285090 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 287058 0 287114 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 289082 0 289138 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 291198 0 291254 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 293222 0 293278 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 295338 0 295394 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 297362 0 297418 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 299386 0 299442 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 301502 0 301558 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 303526 0 303582 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 305550 0 305606 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 307666 0 307722 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 309690 0 309746 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 311806 0 311862 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 313830 0 313886 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 315854 0 315910 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 317970 0 318026 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 319994 0 320050 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 322018 0 322074 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 324134 0 324190 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 326158 0 326214 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 328274 0 328330 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 330298 0 330354 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 332322 0 332378 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 334438 0 334494 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 149150 0 149206 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 161478 0 161534 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 165618 0 165674 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 169758 0 169814 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 173806 0 173862 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 175922 0 175978 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 180062 0 180118 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 182086 0 182142 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 184110 0 184166 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 186226 0 186282 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 188250 0 188306 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 192390 0 192446 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 194414 0 194470 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 198554 0 198610 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 200578 0 200634 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 202694 0 202750 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 206742 0 206798 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 208858 0 208914 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 210882 0 210938 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 212998 0 213054 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 215022 0 215078 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 217046 0 217102 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 219162 0 219218 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 221186 0 221242 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 223210 0 223266 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 225326 0 225382 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 227350 0 227406 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 229466 0 229522 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 231490 0 231546 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 233514 0 233570 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 235630 0 235686 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 237654 0 237710 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 239678 0 239734 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 241794 0 241850 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 243818 0 243874 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 245934 0 245990 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 247958 0 248014 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 249982 0 250038 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 252098 0 252154 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 254122 0 254178 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 256146 0 256202 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 258262 0 258318 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 260286 0 260342 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 262402 0 262458 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 264426 0 264482 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 266450 0 266506 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 268566 0 268622 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 270590 0 270646 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 272614 0 272670 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 274730 0 274786 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 276754 0 276810 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 279514 0 279570 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 281538 0 281594 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 283654 0 283710 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 285678 0 285734 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 287794 0 287850 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 289818 0 289874 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 291842 0 291898 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 293958 0 294014 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 295982 0 296038 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 298006 0 298062 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 94226 0 94282 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 300122 0 300178 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 302146 0 302202 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 304262 0 304318 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 306286 0 306342 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 308310 0 308366 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 310426 0 310482 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 312450 0 312506 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 314474 0 314530 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 316590 0 316646 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 318614 0 318670 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 96342 0 96398 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 320730 0 320786 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 322754 0 322810 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 324778 0 324834 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 326894 0 326950 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 328918 0 328974 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 330942 0 330998 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 333058 0 333114 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 335082 0 335138 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 98366 0 98422 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 100390 0 100446 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 102506 0 102562 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 104530 0 104586 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 108670 0 108726 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 112810 0 112866 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 114834 0 114890 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 116858 0 116914 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 118974 0 119030 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 120998 0 121054 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 127162 0 127218 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 131302 0 131358 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 135442 0 135498 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 137466 0 137522 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 141606 0 141662 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 145746 0 145802 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 147770 0 147826 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 149794 0 149850 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 151910 0 151966 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 156050 0 156106 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 158074 0 158130 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 160098 0 160154 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 162214 0 162270 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 164238 0 164294 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 166262 0 166318 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 168378 0 168434 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 170402 0 170458 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 172518 0 172574 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 174542 0 174598 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 81898 0 81954 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 176566 0 176622 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 178682 0 178738 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 180706 0 180762 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 182730 0 182786 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 184846 0 184902 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 186870 0 186926 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 188986 0 189042 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 191010 0 191066 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 193034 0 193090 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 195150 0 195206 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 197174 0 197230 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 199198 0 199254 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 201314 0 201370 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 203338 0 203394 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 205454 0 205510 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 207478 0 207534 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 209502 0 209558 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 211618 0 211674 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 213642 0 213698 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 215666 0 215722 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 86038 0 86094 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 217782 0 217838 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 219806 0 219862 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 221922 0 221978 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 223946 0 224002 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 225970 0 226026 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 228086 0 228142 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 230110 0 230166 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 232134 0 232190 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 234250 0 234306 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 236274 0 236330 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 238390 0 238446 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 240414 0 240470 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 242438 0 242494 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 244554 0 244610 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 246578 0 246634 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 248602 0 248658 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 250718 0 250774 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 252742 0 252798 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 254858 0 254914 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 256882 0 256938 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 258906 0 258962 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 261022 0 261078 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 263046 0 263102 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 265070 0 265126 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 267186 0 267242 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 269210 0 269266 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 271326 0 271382 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 273350 0 273406 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 275374 0 275430 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 277490 0 277546 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 92202 0 92258 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 74354 0 74410 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 280250 0 280306 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 282274 0 282330 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 284298 0 284354 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 286414 0 286470 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 288438 0 288494 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 290462 0 290518 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 292578 0 292634 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 294602 0 294658 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 296718 0 296774 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 298742 0 298798 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 300766 0 300822 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 302882 0 302938 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 304906 0 304962 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 306930 0 306986 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 309046 0 309102 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 311070 0 311126 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 313186 0 313242 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 315210 0 315266 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 317234 0 317290 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 319350 0 319406 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 321374 0 321430 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 323398 0 323454 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 325514 0 325570 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 327538 0 327594 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 329654 0 329710 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 331678 0 331734 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 333702 0 333758 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 335818 0 335874 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 123758 0 123814 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 136086 0 136142 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 140226 0 140282 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 144366 0 144422 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 148506 0 148562 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 150530 0 150586 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 154670 0 154726 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 164974 0 165030 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 166998 0 167054 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 171138 0 171194 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 177302 0 177358 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 179326 0 179382 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 181442 0 181498 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 183466 0 183522 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 185490 0 185546 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 187606 0 187662 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 189630 0 189686 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 191654 0 191710 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 193770 0 193826 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 195794 0 195850 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 197910 0 197966 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 199934 0 199990 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 201958 0 202014 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 204074 0 204130 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 208122 0 208178 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 210238 0 210294 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 212262 0 212318 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 214378 0 214434 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 216402 0 216458 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 218426 0 218482 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 220542 0 220598 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 222566 0 222622 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 224590 0 224646 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 226706 0 226762 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 228730 0 228786 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 230846 0 230902 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 232870 0 232926 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 234894 0 234950 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 237010 0 237066 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 239034 0 239090 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 241058 0 241114 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 243174 0 243230 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 245198 0 245254 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 247314 0 247370 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 249338 0 249394 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 251362 0 251418 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 253478 0 253534 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 255502 0 255558 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 257526 0 257582 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 259642 0 259698 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 261666 0 261722 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 263782 0 263838 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 265806 0 265862 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 267830 0 267886 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 269946 0 270002 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 271970 0 272026 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 273994 0 274050 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 276110 0 276166 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 278134 0 278190 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 405328 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 405328 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 405328 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 405328 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 405328 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 405328 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 405328 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 405328 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 405328 6 vccd1
port 502 nsew power input
rlabel metal4 s 280688 2128 281008 405328 6 vccd1
port 502 nsew power input
rlabel metal4 s 311408 2128 311728 405328 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 405328 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 405328 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 405328 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 405328 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 405328 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 405328 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 405328 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 405328 6 vssd1
port 503 nsew ground input
rlabel metal4 s 265328 2128 265648 405328 6 vssd1
port 503 nsew ground input
rlabel metal4 s 296048 2128 296368 405328 6 vssd1
port 503 nsew ground input
rlabel metal4 s 326768 2128 327088 405328 6 vssd1
port 503 nsew ground input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 938 0 994 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 72330 0 72386 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 338267 407623
string LEFview TRUE
string GDS_FILE /project/openlane/user_project/runs/user_project/results/magic/user_project.gds
string GDS_END 157956112
string GDS_START 1045048
<< end >>

