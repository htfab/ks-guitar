VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project
  CLASS BLOCK ;
  FOREIGN user_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 1691.335 BY 2038.115 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 2034.115 7.730 2038.115 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 2034.115 452.550 2038.115 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 2034.115 497.170 2038.115 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 2034.115 541.790 2038.115 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 2034.115 585.950 2038.115 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 2034.115 630.570 2038.115 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 2034.115 675.190 2038.115 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 2034.115 719.810 2038.115 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 2034.115 763.970 2038.115 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 2034.115 808.590 2038.115 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.930 2034.115 853.210 2038.115 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 2034.115 51.890 2038.115 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 2034.115 897.830 2038.115 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 2034.115 942.450 2038.115 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.330 2034.115 986.610 2038.115 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.950 2034.115 1031.230 2038.115 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.570 2034.115 1075.850 2038.115 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.190 2034.115 1120.470 2038.115 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.350 2034.115 1164.630 2038.115 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.970 2034.115 1209.250 2038.115 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.590 2034.115 1253.870 2038.115 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.210 2034.115 1298.490 2038.115 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 2034.115 96.510 2038.115 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.370 2034.115 1342.650 2038.115 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.990 2034.115 1387.270 2038.115 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.610 2034.115 1431.890 2038.115 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.230 2034.115 1476.510 2038.115 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1520.390 2034.115 1520.670 2038.115 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.010 2034.115 1565.290 2038.115 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1609.630 2034.115 1609.910 2038.115 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.250 2034.115 1654.530 2038.115 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 2034.115 141.130 2038.115 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 2034.115 185.750 2038.115 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 2034.115 229.910 2038.115 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 2034.115 274.530 2038.115 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 2034.115 319.150 2038.115 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 2034.115 363.770 2038.115 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 2034.115 407.930 2038.115 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 2034.115 22.450 2038.115 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 2034.115 467.270 2038.115 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 2034.115 511.890 2038.115 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 2034.115 556.510 2038.115 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 2034.115 601.130 2038.115 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 2034.115 645.290 2038.115 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 2034.115 689.910 2038.115 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 2034.115 734.530 2038.115 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 2034.115 779.150 2038.115 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.030 2034.115 823.310 2038.115 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.650 2034.115 867.930 2038.115 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 2034.115 67.070 2038.115 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.270 2034.115 912.550 2038.115 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.890 2034.115 957.170 2038.115 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 2034.115 1001.790 2038.115 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.670 2034.115 1045.950 2038.115 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.290 2034.115 1090.570 2038.115 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.910 2034.115 1135.190 2038.115 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.530 2034.115 1179.810 2038.115 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 2034.115 1223.970 2038.115 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.310 2034.115 1268.590 2038.115 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.930 2034.115 1313.210 2038.115 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 2034.115 111.230 2038.115 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.550 2034.115 1357.830 2038.115 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.710 2034.115 1401.990 2038.115 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.330 2034.115 1446.610 2038.115 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 2034.115 1491.230 2038.115 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.570 2034.115 1535.850 2038.115 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.730 2034.115 1580.010 2038.115 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1624.350 2034.115 1624.630 2038.115 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.970 2034.115 1669.250 2038.115 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 2034.115 155.850 2038.115 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 2034.115 200.470 2038.115 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 2034.115 245.090 2038.115 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 2034.115 289.250 2038.115 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 2034.115 333.870 2038.115 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 2034.115 378.490 2038.115 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 2034.115 423.110 2038.115 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 2034.115 37.170 2038.115 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 2034.115 482.450 2038.115 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 2034.115 526.610 2038.115 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 2034.115 571.230 2038.115 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 2034.115 615.850 2038.115 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 2034.115 660.470 2038.115 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 2034.115 704.630 2038.115 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 2034.115 749.250 2038.115 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 2034.115 793.870 2038.115 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 2034.115 838.490 2038.115 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.830 2034.115 883.110 2038.115 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 2034.115 81.790 2038.115 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.990 2034.115 927.270 2038.115 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.610 2034.115 971.890 2038.115 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.230 2034.115 1016.510 2038.115 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.850 2034.115 1061.130 2038.115 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.010 2034.115 1105.290 2038.115 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 2034.115 1149.910 2038.115 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.250 2034.115 1194.530 2038.115 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.870 2034.115 1239.150 2038.115 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.030 2034.115 1283.310 2038.115 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.650 2034.115 1327.930 2038.115 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 2034.115 126.410 2038.115 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1372.270 2034.115 1372.550 2038.115 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 2034.115 1417.170 2038.115 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.050 2034.115 1461.330 2038.115 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1505.670 2034.115 1505.950 2038.115 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.290 2034.115 1550.570 2038.115 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.910 2034.115 1595.190 2038.115 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.070 2034.115 1639.350 2038.115 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.690 2034.115 1683.970 2038.115 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 2034.115 170.570 2038.115 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 2034.115 215.190 2038.115 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 2034.115 259.810 2038.115 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 2034.115 304.430 2038.115 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 2034.115 348.590 2038.115 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 2034.115 393.210 2038.115 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 2034.115 437.830 2038.115 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1682.310 0.000 1682.590 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.990 0.000 1686.270 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.210 0.000 1689.490 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 0.000 365.150 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.350 0.000 1394.630 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.470 0.000 1404.750 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.590 0.000 1414.870 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1425.170 0.000 1425.450 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.290 0.000 1435.570 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.410 0.000 1445.690 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.990 0.000 1456.270 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1466.110 0.000 1466.390 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.690 0.000 1476.970 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.810 0.000 1487.090 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.930 0.000 1497.210 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.510 0.000 1507.790 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.630 0.000 1517.910 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.750 0.000 1528.030 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1538.330 0.000 1538.610 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.450 0.000 1548.730 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.030 0.000 1559.310 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.150 0.000 1569.430 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.270 0.000 1579.550 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.850 0.000 1590.130 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 0.000 478.310 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.970 0.000 1600.250 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.090 0.000 1610.370 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.670 0.000 1620.950 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1630.790 0.000 1631.070 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1641.370 0.000 1641.650 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.490 0.000 1651.770 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.610 0.000 1661.890 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.190 0.000 1672.470 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 0.000 499.010 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 0.000 550.530 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 0.000 571.230 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 0.000 602.050 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 0.000 622.290 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 0.000 632.870 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 0.000 642.990 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 0.000 673.810 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 0.000 684.390 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 0.000 704.630 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 0.000 725.330 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 0.000 735.910 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 0.000 746.030 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.870 0.000 756.150 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 0.000 776.850 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 0.000 786.970 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 0.000 797.550 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 0.000 807.670 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 0.000 828.370 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 0.000 838.490 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 0.000 849.070 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.910 0.000 859.190 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.030 0.000 869.310 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 0.000 879.890 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.730 0.000 890.010 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.310 0.000 900.590 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.430 0.000 910.710 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 0.000 920.830 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 0.000 931.410 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.250 0.000 941.530 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.370 0.000 951.650 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.950 0.000 962.230 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.070 0.000 972.350 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 0.000 982.930 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.770 0.000 993.050 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.890 0.000 1003.170 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.470 0.000 1013.750 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.590 0.000 1023.870 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.290 0.000 1044.570 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.410 0.000 1054.690 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.990 0.000 1065.270 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.110 0.000 1075.390 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 0.000 1085.510 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.810 0.000 1096.090 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.930 0.000 1106.210 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.050 0.000 1116.330 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.630 0.000 1126.910 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 0.000 1137.030 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.330 0.000 1147.610 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.450 0.000 1157.730 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.570 0.000 1167.850 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.150 0.000 1178.430 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 0.000 1188.550 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.390 0.000 1198.670 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.970 0.000 1209.250 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.090 0.000 1219.370 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.670 0.000 1229.950 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 0.000 1240.070 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.910 0.000 1250.190 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.490 0.000 1260.770 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1270.610 0.000 1270.890 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.730 0.000 1281.010 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.430 0.000 1301.710 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.010 0.000 1312.290 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.130 0.000 1322.410 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.250 0.000 1332.530 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 0.000 1343.110 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.950 0.000 1353.230 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.070 0.000 1363.350 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.650 0.000 1373.930 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1383.770 0.000 1384.050 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 0.000 1397.850 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.690 0.000 1407.970 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.270 0.000 1418.550 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.390 0.000 1428.670 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.970 0.000 1439.250 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 0.000 1449.370 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.210 0.000 1459.490 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1469.790 0.000 1470.070 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.910 0.000 1480.190 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.030 0.000 1490.310 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.610 0.000 1500.890 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.730 0.000 1511.010 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.310 0.000 1521.590 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1531.430 0.000 1531.710 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1541.550 0.000 1541.830 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.130 0.000 1552.410 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.250 0.000 1562.530 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.370 0.000 1572.650 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1582.950 0.000 1583.230 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.070 0.000 1593.350 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.650 0.000 1603.930 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.770 0.000 1614.050 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1623.890 0.000 1624.170 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.470 0.000 1634.750 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.590 0.000 1644.870 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.710 0.000 1654.990 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1665.290 0.000 1665.570 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.410 0.000 1675.690 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 0.000 492.110 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 0.000 533.510 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 0.000 543.630 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 0.000 564.330 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 0.000 584.570 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 0.000 595.150 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 0.000 605.270 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 0.000 625.970 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 0.000 646.670 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 0.000 677.490 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 0.000 687.610 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 0.000 698.190 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 0.000 708.310 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 0.000 729.010 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 0.000 739.130 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 0.000 749.250 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.550 0.000 759.830 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 0.000 780.530 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.370 0.000 790.650 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 0.000 800.770 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 0.000 811.350 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 0.000 831.590 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 0.000 842.170 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.010 0.000 852.290 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 0.000 862.870 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 0.000 872.990 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.830 0.000 883.110 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 0.000 893.690 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.530 0.000 903.810 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 0.000 913.930 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 0.000 924.510 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.350 0.000 934.630 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.930 0.000 945.210 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 0.000 955.330 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.170 0.000 965.450 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.870 0.000 986.150 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.990 0.000 996.270 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.570 0.000 1006.850 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.690 0.000 1016.970 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 0.000 1027.550 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 0.000 1037.670 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.510 0.000 1047.790 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.090 0.000 1058.370 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.210 0.000 1068.490 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.330 0.000 1078.610 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.910 0.000 1089.190 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.030 0.000 1099.310 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.610 0.000 1109.890 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.730 0.000 1120.010 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1129.850 0.000 1130.130 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.430 0.000 1140.710 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.550 0.000 1150.830 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.670 0.000 1160.950 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.250 0.000 1171.530 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.370 0.000 1181.650 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.950 0.000 1192.230 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.070 0.000 1202.350 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1212.190 0.000 1212.470 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1222.770 0.000 1223.050 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.890 0.000 1233.170 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.010 0.000 1243.290 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.590 0.000 1253.870 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.710 0.000 1263.990 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.290 0.000 1274.570 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.410 0.000 1284.690 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 0.000 1294.810 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.110 0.000 1305.390 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.230 0.000 1315.510 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1325.350 0.000 1325.630 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.930 0.000 1336.210 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 0.000 1346.330 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.630 0.000 1356.910 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.750 0.000 1367.030 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.870 0.000 1377.150 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.450 0.000 1387.730 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.250 0.000 1401.530 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1411.370 0.000 1411.650 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.490 0.000 1421.770 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.070 0.000 1432.350 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.190 0.000 1442.470 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 0.000 1452.590 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.890 0.000 1463.170 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.010 0.000 1473.290 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.590 0.000 1483.870 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1493.710 0.000 1493.990 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.830 0.000 1504.110 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.410 0.000 1514.690 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.530 0.000 1524.810 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.650 0.000 1534.930 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.230 0.000 1545.510 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 0.000 1555.630 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.930 0.000 1566.210 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.050 0.000 1576.330 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.170 0.000 1586.450 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.750 0.000 1597.030 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.870 0.000 1607.150 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.990 0.000 1617.270 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.570 0.000 1627.850 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1637.690 0.000 1637.970 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.270 0.000 1648.550 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.390 0.000 1658.670 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.510 0.000 1668.790 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.090 0.000 1679.370 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 0.000 526.610 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 0.000 546.850 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 0.000 567.550 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 0.000 619.070 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 0.000 629.190 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 0.000 639.770 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 0.000 670.590 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 0.000 701.410 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 0.000 711.530 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 0.000 722.110 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.950 0.000 732.230 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 0.000 742.810 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 0.000 752.930 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 0.000 763.050 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 0.000 773.630 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.470 0.000 783.750 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.170 0.000 804.450 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 0.000 814.570 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.870 0.000 825.150 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.990 0.000 835.270 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.110 0.000 845.390 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 0.000 855.970 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 0.000 866.090 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 0.000 876.210 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.510 0.000 886.790 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.630 0.000 896.910 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.210 0.000 907.490 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.330 0.000 917.610 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.030 0.000 938.310 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.150 0.000 948.430 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.270 0.000 958.550 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.850 0.000 969.130 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.550 0.000 989.830 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.670 0.000 999.950 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.790 0.000 1010.070 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.370 0.000 1020.650 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 0.000 1030.770 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.610 0.000 1040.890 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.190 0.000 1051.470 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.310 0.000 1061.590 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.890 0.000 1072.170 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.130 0.000 1092.410 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.710 0.000 1102.990 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.830 0.000 1113.110 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.950 0.000 1123.230 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.530 0.000 1133.810 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.650 0.000 1143.930 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.230 0.000 1154.510 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.350 0.000 1164.630 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.470 0.000 1174.750 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 0.000 1185.330 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.170 0.000 1195.450 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.290 0.000 1205.570 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.870 0.000 1216.150 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.990 0.000 1226.270 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.570 0.000 1236.850 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.690 0.000 1246.970 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.810 0.000 1257.090 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.390 0.000 1267.670 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.510 0.000 1277.790 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.630 0.000 1287.910 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.210 0.000 1298.490 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.330 0.000 1308.610 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.910 0.000 1319.190 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.030 0.000 1329.310 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.150 0.000 1339.430 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.730 0.000 1350.010 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.850 0.000 1360.130 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.970 0.000 1370.250 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.550 0.000 1380.830 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.670 0.000 1390.950 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 0.000 464.510 4.000 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 2026.640 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 2026.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 2026.640 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 1685.440 2026.485 ;
      LAYER met1 ;
        RECT 1.450 6.840 1689.510 2028.400 ;
      LAYER met2 ;
        RECT 1.480 2033.835 7.170 2034.290 ;
        RECT 8.010 2033.835 21.890 2034.290 ;
        RECT 22.730 2033.835 36.610 2034.290 ;
        RECT 37.450 2033.835 51.330 2034.290 ;
        RECT 52.170 2033.835 66.510 2034.290 ;
        RECT 67.350 2033.835 81.230 2034.290 ;
        RECT 82.070 2033.835 95.950 2034.290 ;
        RECT 96.790 2033.835 110.670 2034.290 ;
        RECT 111.510 2033.835 125.850 2034.290 ;
        RECT 126.690 2033.835 140.570 2034.290 ;
        RECT 141.410 2033.835 155.290 2034.290 ;
        RECT 156.130 2033.835 170.010 2034.290 ;
        RECT 170.850 2033.835 185.190 2034.290 ;
        RECT 186.030 2033.835 199.910 2034.290 ;
        RECT 200.750 2033.835 214.630 2034.290 ;
        RECT 215.470 2033.835 229.350 2034.290 ;
        RECT 230.190 2033.835 244.530 2034.290 ;
        RECT 245.370 2033.835 259.250 2034.290 ;
        RECT 260.090 2033.835 273.970 2034.290 ;
        RECT 274.810 2033.835 288.690 2034.290 ;
        RECT 289.530 2033.835 303.870 2034.290 ;
        RECT 304.710 2033.835 318.590 2034.290 ;
        RECT 319.430 2033.835 333.310 2034.290 ;
        RECT 334.150 2033.835 348.030 2034.290 ;
        RECT 348.870 2033.835 363.210 2034.290 ;
        RECT 364.050 2033.835 377.930 2034.290 ;
        RECT 378.770 2033.835 392.650 2034.290 ;
        RECT 393.490 2033.835 407.370 2034.290 ;
        RECT 408.210 2033.835 422.550 2034.290 ;
        RECT 423.390 2033.835 437.270 2034.290 ;
        RECT 438.110 2033.835 451.990 2034.290 ;
        RECT 452.830 2033.835 466.710 2034.290 ;
        RECT 467.550 2033.835 481.890 2034.290 ;
        RECT 482.730 2033.835 496.610 2034.290 ;
        RECT 497.450 2033.835 511.330 2034.290 ;
        RECT 512.170 2033.835 526.050 2034.290 ;
        RECT 526.890 2033.835 541.230 2034.290 ;
        RECT 542.070 2033.835 555.950 2034.290 ;
        RECT 556.790 2033.835 570.670 2034.290 ;
        RECT 571.510 2033.835 585.390 2034.290 ;
        RECT 586.230 2033.835 600.570 2034.290 ;
        RECT 601.410 2033.835 615.290 2034.290 ;
        RECT 616.130 2033.835 630.010 2034.290 ;
        RECT 630.850 2033.835 644.730 2034.290 ;
        RECT 645.570 2033.835 659.910 2034.290 ;
        RECT 660.750 2033.835 674.630 2034.290 ;
        RECT 675.470 2033.835 689.350 2034.290 ;
        RECT 690.190 2033.835 704.070 2034.290 ;
        RECT 704.910 2033.835 719.250 2034.290 ;
        RECT 720.090 2033.835 733.970 2034.290 ;
        RECT 734.810 2033.835 748.690 2034.290 ;
        RECT 749.530 2033.835 763.410 2034.290 ;
        RECT 764.250 2033.835 778.590 2034.290 ;
        RECT 779.430 2033.835 793.310 2034.290 ;
        RECT 794.150 2033.835 808.030 2034.290 ;
        RECT 808.870 2033.835 822.750 2034.290 ;
        RECT 823.590 2033.835 837.930 2034.290 ;
        RECT 838.770 2033.835 852.650 2034.290 ;
        RECT 853.490 2033.835 867.370 2034.290 ;
        RECT 868.210 2033.835 882.550 2034.290 ;
        RECT 883.390 2033.835 897.270 2034.290 ;
        RECT 898.110 2033.835 911.990 2034.290 ;
        RECT 912.830 2033.835 926.710 2034.290 ;
        RECT 927.550 2033.835 941.890 2034.290 ;
        RECT 942.730 2033.835 956.610 2034.290 ;
        RECT 957.450 2033.835 971.330 2034.290 ;
        RECT 972.170 2033.835 986.050 2034.290 ;
        RECT 986.890 2033.835 1001.230 2034.290 ;
        RECT 1002.070 2033.835 1015.950 2034.290 ;
        RECT 1016.790 2033.835 1030.670 2034.290 ;
        RECT 1031.510 2033.835 1045.390 2034.290 ;
        RECT 1046.230 2033.835 1060.570 2034.290 ;
        RECT 1061.410 2033.835 1075.290 2034.290 ;
        RECT 1076.130 2033.835 1090.010 2034.290 ;
        RECT 1090.850 2033.835 1104.730 2034.290 ;
        RECT 1105.570 2033.835 1119.910 2034.290 ;
        RECT 1120.750 2033.835 1134.630 2034.290 ;
        RECT 1135.470 2033.835 1149.350 2034.290 ;
        RECT 1150.190 2033.835 1164.070 2034.290 ;
        RECT 1164.910 2033.835 1179.250 2034.290 ;
        RECT 1180.090 2033.835 1193.970 2034.290 ;
        RECT 1194.810 2033.835 1208.690 2034.290 ;
        RECT 1209.530 2033.835 1223.410 2034.290 ;
        RECT 1224.250 2033.835 1238.590 2034.290 ;
        RECT 1239.430 2033.835 1253.310 2034.290 ;
        RECT 1254.150 2033.835 1268.030 2034.290 ;
        RECT 1268.870 2033.835 1282.750 2034.290 ;
        RECT 1283.590 2033.835 1297.930 2034.290 ;
        RECT 1298.770 2033.835 1312.650 2034.290 ;
        RECT 1313.490 2033.835 1327.370 2034.290 ;
        RECT 1328.210 2033.835 1342.090 2034.290 ;
        RECT 1342.930 2033.835 1357.270 2034.290 ;
        RECT 1358.110 2033.835 1371.990 2034.290 ;
        RECT 1372.830 2033.835 1386.710 2034.290 ;
        RECT 1387.550 2033.835 1401.430 2034.290 ;
        RECT 1402.270 2033.835 1416.610 2034.290 ;
        RECT 1417.450 2033.835 1431.330 2034.290 ;
        RECT 1432.170 2033.835 1446.050 2034.290 ;
        RECT 1446.890 2033.835 1460.770 2034.290 ;
        RECT 1461.610 2033.835 1475.950 2034.290 ;
        RECT 1476.790 2033.835 1490.670 2034.290 ;
        RECT 1491.510 2033.835 1505.390 2034.290 ;
        RECT 1506.230 2033.835 1520.110 2034.290 ;
        RECT 1520.950 2033.835 1535.290 2034.290 ;
        RECT 1536.130 2033.835 1550.010 2034.290 ;
        RECT 1550.850 2033.835 1564.730 2034.290 ;
        RECT 1565.570 2033.835 1579.450 2034.290 ;
        RECT 1580.290 2033.835 1594.630 2034.290 ;
        RECT 1595.470 2033.835 1609.350 2034.290 ;
        RECT 1610.190 2033.835 1624.070 2034.290 ;
        RECT 1624.910 2033.835 1638.790 2034.290 ;
        RECT 1639.630 2033.835 1653.970 2034.290 ;
        RECT 1654.810 2033.835 1668.690 2034.290 ;
        RECT 1669.530 2033.835 1683.410 2034.290 ;
        RECT 1684.250 2033.835 1689.480 2034.290 ;
        RECT 1.480 4.280 1689.480 2033.835 ;
        RECT 2.030 3.670 4.410 4.280 ;
        RECT 5.250 3.670 7.630 4.280 ;
        RECT 8.470 3.670 11.310 4.280 ;
        RECT 12.150 3.670 14.530 4.280 ;
        RECT 15.370 3.670 18.210 4.280 ;
        RECT 19.050 3.670 21.430 4.280 ;
        RECT 22.270 3.670 25.110 4.280 ;
        RECT 25.950 3.670 28.330 4.280 ;
        RECT 29.170 3.670 32.010 4.280 ;
        RECT 32.850 3.670 35.230 4.280 ;
        RECT 36.070 3.670 38.910 4.280 ;
        RECT 39.750 3.670 42.130 4.280 ;
        RECT 42.970 3.670 45.350 4.280 ;
        RECT 46.190 3.670 49.030 4.280 ;
        RECT 49.870 3.670 52.250 4.280 ;
        RECT 53.090 3.670 55.930 4.280 ;
        RECT 56.770 3.670 59.150 4.280 ;
        RECT 59.990 3.670 62.830 4.280 ;
        RECT 63.670 3.670 66.050 4.280 ;
        RECT 66.890 3.670 69.730 4.280 ;
        RECT 70.570 3.670 72.950 4.280 ;
        RECT 73.790 3.670 76.630 4.280 ;
        RECT 77.470 3.670 79.850 4.280 ;
        RECT 80.690 3.670 83.530 4.280 ;
        RECT 84.370 3.670 86.750 4.280 ;
        RECT 87.590 3.670 89.970 4.280 ;
        RECT 90.810 3.670 93.650 4.280 ;
        RECT 94.490 3.670 96.870 4.280 ;
        RECT 97.710 3.670 100.550 4.280 ;
        RECT 101.390 3.670 103.770 4.280 ;
        RECT 104.610 3.670 107.450 4.280 ;
        RECT 108.290 3.670 110.670 4.280 ;
        RECT 111.510 3.670 114.350 4.280 ;
        RECT 115.190 3.670 117.570 4.280 ;
        RECT 118.410 3.670 121.250 4.280 ;
        RECT 122.090 3.670 124.470 4.280 ;
        RECT 125.310 3.670 127.690 4.280 ;
        RECT 128.530 3.670 131.370 4.280 ;
        RECT 132.210 3.670 134.590 4.280 ;
        RECT 135.430 3.670 138.270 4.280 ;
        RECT 139.110 3.670 141.490 4.280 ;
        RECT 142.330 3.670 145.170 4.280 ;
        RECT 146.010 3.670 148.390 4.280 ;
        RECT 149.230 3.670 152.070 4.280 ;
        RECT 152.910 3.670 155.290 4.280 ;
        RECT 156.130 3.670 158.970 4.280 ;
        RECT 159.810 3.670 162.190 4.280 ;
        RECT 163.030 3.670 165.870 4.280 ;
        RECT 166.710 3.670 169.090 4.280 ;
        RECT 169.930 3.670 172.310 4.280 ;
        RECT 173.150 3.670 175.990 4.280 ;
        RECT 176.830 3.670 179.210 4.280 ;
        RECT 180.050 3.670 182.890 4.280 ;
        RECT 183.730 3.670 186.110 4.280 ;
        RECT 186.950 3.670 189.790 4.280 ;
        RECT 190.630 3.670 193.010 4.280 ;
        RECT 193.850 3.670 196.690 4.280 ;
        RECT 197.530 3.670 199.910 4.280 ;
        RECT 200.750 3.670 203.590 4.280 ;
        RECT 204.430 3.670 206.810 4.280 ;
        RECT 207.650 3.670 210.030 4.280 ;
        RECT 210.870 3.670 213.710 4.280 ;
        RECT 214.550 3.670 216.930 4.280 ;
        RECT 217.770 3.670 220.610 4.280 ;
        RECT 221.450 3.670 223.830 4.280 ;
        RECT 224.670 3.670 227.510 4.280 ;
        RECT 228.350 3.670 230.730 4.280 ;
        RECT 231.570 3.670 234.410 4.280 ;
        RECT 235.250 3.670 237.630 4.280 ;
        RECT 238.470 3.670 241.310 4.280 ;
        RECT 242.150 3.670 244.530 4.280 ;
        RECT 245.370 3.670 248.210 4.280 ;
        RECT 249.050 3.670 251.430 4.280 ;
        RECT 252.270 3.670 254.650 4.280 ;
        RECT 255.490 3.670 258.330 4.280 ;
        RECT 259.170 3.670 261.550 4.280 ;
        RECT 262.390 3.670 265.230 4.280 ;
        RECT 266.070 3.670 268.450 4.280 ;
        RECT 269.290 3.670 272.130 4.280 ;
        RECT 272.970 3.670 275.350 4.280 ;
        RECT 276.190 3.670 279.030 4.280 ;
        RECT 279.870 3.670 282.250 4.280 ;
        RECT 283.090 3.670 285.930 4.280 ;
        RECT 286.770 3.670 289.150 4.280 ;
        RECT 289.990 3.670 292.370 4.280 ;
        RECT 293.210 3.670 296.050 4.280 ;
        RECT 296.890 3.670 299.270 4.280 ;
        RECT 300.110 3.670 302.950 4.280 ;
        RECT 303.790 3.670 306.170 4.280 ;
        RECT 307.010 3.670 309.850 4.280 ;
        RECT 310.690 3.670 313.070 4.280 ;
        RECT 313.910 3.670 316.750 4.280 ;
        RECT 317.590 3.670 319.970 4.280 ;
        RECT 320.810 3.670 323.650 4.280 ;
        RECT 324.490 3.670 326.870 4.280 ;
        RECT 327.710 3.670 330.550 4.280 ;
        RECT 331.390 3.670 333.770 4.280 ;
        RECT 334.610 3.670 336.990 4.280 ;
        RECT 337.830 3.670 340.670 4.280 ;
        RECT 341.510 3.670 343.890 4.280 ;
        RECT 344.730 3.670 347.570 4.280 ;
        RECT 348.410 3.670 350.790 4.280 ;
        RECT 351.630 3.670 354.470 4.280 ;
        RECT 355.310 3.670 357.690 4.280 ;
        RECT 358.530 3.670 361.370 4.280 ;
        RECT 362.210 3.670 364.590 4.280 ;
        RECT 365.430 3.670 368.270 4.280 ;
        RECT 369.110 3.670 371.490 4.280 ;
        RECT 372.330 3.670 374.710 4.280 ;
        RECT 375.550 3.670 378.390 4.280 ;
        RECT 379.230 3.670 381.610 4.280 ;
        RECT 382.450 3.670 385.290 4.280 ;
        RECT 386.130 3.670 388.510 4.280 ;
        RECT 389.350 3.670 392.190 4.280 ;
        RECT 393.030 3.670 395.410 4.280 ;
        RECT 396.250 3.670 399.090 4.280 ;
        RECT 399.930 3.670 402.310 4.280 ;
        RECT 403.150 3.670 405.990 4.280 ;
        RECT 406.830 3.670 409.210 4.280 ;
        RECT 410.050 3.670 412.890 4.280 ;
        RECT 413.730 3.670 416.110 4.280 ;
        RECT 416.950 3.670 419.330 4.280 ;
        RECT 420.170 3.670 423.010 4.280 ;
        RECT 423.850 3.670 426.230 4.280 ;
        RECT 427.070 3.670 429.910 4.280 ;
        RECT 430.750 3.670 433.130 4.280 ;
        RECT 433.970 3.670 436.810 4.280 ;
        RECT 437.650 3.670 440.030 4.280 ;
        RECT 440.870 3.670 443.710 4.280 ;
        RECT 444.550 3.670 446.930 4.280 ;
        RECT 447.770 3.670 450.610 4.280 ;
        RECT 451.450 3.670 453.830 4.280 ;
        RECT 454.670 3.670 457.050 4.280 ;
        RECT 457.890 3.670 460.730 4.280 ;
        RECT 461.570 3.670 463.950 4.280 ;
        RECT 464.790 3.670 467.630 4.280 ;
        RECT 468.470 3.670 470.850 4.280 ;
        RECT 471.690 3.670 474.530 4.280 ;
        RECT 475.370 3.670 477.750 4.280 ;
        RECT 478.590 3.670 481.430 4.280 ;
        RECT 482.270 3.670 484.650 4.280 ;
        RECT 485.490 3.670 488.330 4.280 ;
        RECT 489.170 3.670 491.550 4.280 ;
        RECT 492.390 3.670 495.230 4.280 ;
        RECT 496.070 3.670 498.450 4.280 ;
        RECT 499.290 3.670 501.670 4.280 ;
        RECT 502.510 3.670 505.350 4.280 ;
        RECT 506.190 3.670 508.570 4.280 ;
        RECT 509.410 3.670 512.250 4.280 ;
        RECT 513.090 3.670 515.470 4.280 ;
        RECT 516.310 3.670 519.150 4.280 ;
        RECT 519.990 3.670 522.370 4.280 ;
        RECT 523.210 3.670 526.050 4.280 ;
        RECT 526.890 3.670 529.270 4.280 ;
        RECT 530.110 3.670 532.950 4.280 ;
        RECT 533.790 3.670 536.170 4.280 ;
        RECT 537.010 3.670 539.390 4.280 ;
        RECT 540.230 3.670 543.070 4.280 ;
        RECT 543.910 3.670 546.290 4.280 ;
        RECT 547.130 3.670 549.970 4.280 ;
        RECT 550.810 3.670 553.190 4.280 ;
        RECT 554.030 3.670 556.870 4.280 ;
        RECT 557.710 3.670 560.090 4.280 ;
        RECT 560.930 3.670 563.770 4.280 ;
        RECT 564.610 3.670 566.990 4.280 ;
        RECT 567.830 3.670 570.670 4.280 ;
        RECT 571.510 3.670 573.890 4.280 ;
        RECT 574.730 3.670 577.570 4.280 ;
        RECT 578.410 3.670 580.790 4.280 ;
        RECT 581.630 3.670 584.010 4.280 ;
        RECT 584.850 3.670 587.690 4.280 ;
        RECT 588.530 3.670 590.910 4.280 ;
        RECT 591.750 3.670 594.590 4.280 ;
        RECT 595.430 3.670 597.810 4.280 ;
        RECT 598.650 3.670 601.490 4.280 ;
        RECT 602.330 3.670 604.710 4.280 ;
        RECT 605.550 3.670 608.390 4.280 ;
        RECT 609.230 3.670 611.610 4.280 ;
        RECT 612.450 3.670 615.290 4.280 ;
        RECT 616.130 3.670 618.510 4.280 ;
        RECT 619.350 3.670 621.730 4.280 ;
        RECT 622.570 3.670 625.410 4.280 ;
        RECT 626.250 3.670 628.630 4.280 ;
        RECT 629.470 3.670 632.310 4.280 ;
        RECT 633.150 3.670 635.530 4.280 ;
        RECT 636.370 3.670 639.210 4.280 ;
        RECT 640.050 3.670 642.430 4.280 ;
        RECT 643.270 3.670 646.110 4.280 ;
        RECT 646.950 3.670 649.330 4.280 ;
        RECT 650.170 3.670 653.010 4.280 ;
        RECT 653.850 3.670 656.230 4.280 ;
        RECT 657.070 3.670 659.910 4.280 ;
        RECT 660.750 3.670 663.130 4.280 ;
        RECT 663.970 3.670 666.350 4.280 ;
        RECT 667.190 3.670 670.030 4.280 ;
        RECT 670.870 3.670 673.250 4.280 ;
        RECT 674.090 3.670 676.930 4.280 ;
        RECT 677.770 3.670 680.150 4.280 ;
        RECT 680.990 3.670 683.830 4.280 ;
        RECT 684.670 3.670 687.050 4.280 ;
        RECT 687.890 3.670 690.730 4.280 ;
        RECT 691.570 3.670 693.950 4.280 ;
        RECT 694.790 3.670 697.630 4.280 ;
        RECT 698.470 3.670 700.850 4.280 ;
        RECT 701.690 3.670 704.070 4.280 ;
        RECT 704.910 3.670 707.750 4.280 ;
        RECT 708.590 3.670 710.970 4.280 ;
        RECT 711.810 3.670 714.650 4.280 ;
        RECT 715.490 3.670 717.870 4.280 ;
        RECT 718.710 3.670 721.550 4.280 ;
        RECT 722.390 3.670 724.770 4.280 ;
        RECT 725.610 3.670 728.450 4.280 ;
        RECT 729.290 3.670 731.670 4.280 ;
        RECT 732.510 3.670 735.350 4.280 ;
        RECT 736.190 3.670 738.570 4.280 ;
        RECT 739.410 3.670 742.250 4.280 ;
        RECT 743.090 3.670 745.470 4.280 ;
        RECT 746.310 3.670 748.690 4.280 ;
        RECT 749.530 3.670 752.370 4.280 ;
        RECT 753.210 3.670 755.590 4.280 ;
        RECT 756.430 3.670 759.270 4.280 ;
        RECT 760.110 3.670 762.490 4.280 ;
        RECT 763.330 3.670 766.170 4.280 ;
        RECT 767.010 3.670 769.390 4.280 ;
        RECT 770.230 3.670 773.070 4.280 ;
        RECT 773.910 3.670 776.290 4.280 ;
        RECT 777.130 3.670 779.970 4.280 ;
        RECT 780.810 3.670 783.190 4.280 ;
        RECT 784.030 3.670 786.410 4.280 ;
        RECT 787.250 3.670 790.090 4.280 ;
        RECT 790.930 3.670 793.310 4.280 ;
        RECT 794.150 3.670 796.990 4.280 ;
        RECT 797.830 3.670 800.210 4.280 ;
        RECT 801.050 3.670 803.890 4.280 ;
        RECT 804.730 3.670 807.110 4.280 ;
        RECT 807.950 3.670 810.790 4.280 ;
        RECT 811.630 3.670 814.010 4.280 ;
        RECT 814.850 3.670 817.690 4.280 ;
        RECT 818.530 3.670 820.910 4.280 ;
        RECT 821.750 3.670 824.590 4.280 ;
        RECT 825.430 3.670 827.810 4.280 ;
        RECT 828.650 3.670 831.030 4.280 ;
        RECT 831.870 3.670 834.710 4.280 ;
        RECT 835.550 3.670 837.930 4.280 ;
        RECT 838.770 3.670 841.610 4.280 ;
        RECT 842.450 3.670 844.830 4.280 ;
        RECT 845.670 3.670 848.510 4.280 ;
        RECT 849.350 3.670 851.730 4.280 ;
        RECT 852.570 3.670 855.410 4.280 ;
        RECT 856.250 3.670 858.630 4.280 ;
        RECT 859.470 3.670 862.310 4.280 ;
        RECT 863.150 3.670 865.530 4.280 ;
        RECT 866.370 3.670 868.750 4.280 ;
        RECT 869.590 3.670 872.430 4.280 ;
        RECT 873.270 3.670 875.650 4.280 ;
        RECT 876.490 3.670 879.330 4.280 ;
        RECT 880.170 3.670 882.550 4.280 ;
        RECT 883.390 3.670 886.230 4.280 ;
        RECT 887.070 3.670 889.450 4.280 ;
        RECT 890.290 3.670 893.130 4.280 ;
        RECT 893.970 3.670 896.350 4.280 ;
        RECT 897.190 3.670 900.030 4.280 ;
        RECT 900.870 3.670 903.250 4.280 ;
        RECT 904.090 3.670 906.930 4.280 ;
        RECT 907.770 3.670 910.150 4.280 ;
        RECT 910.990 3.670 913.370 4.280 ;
        RECT 914.210 3.670 917.050 4.280 ;
        RECT 917.890 3.670 920.270 4.280 ;
        RECT 921.110 3.670 923.950 4.280 ;
        RECT 924.790 3.670 927.170 4.280 ;
        RECT 928.010 3.670 930.850 4.280 ;
        RECT 931.690 3.670 934.070 4.280 ;
        RECT 934.910 3.670 937.750 4.280 ;
        RECT 938.590 3.670 940.970 4.280 ;
        RECT 941.810 3.670 944.650 4.280 ;
        RECT 945.490 3.670 947.870 4.280 ;
        RECT 948.710 3.670 951.090 4.280 ;
        RECT 951.930 3.670 954.770 4.280 ;
        RECT 955.610 3.670 957.990 4.280 ;
        RECT 958.830 3.670 961.670 4.280 ;
        RECT 962.510 3.670 964.890 4.280 ;
        RECT 965.730 3.670 968.570 4.280 ;
        RECT 969.410 3.670 971.790 4.280 ;
        RECT 972.630 3.670 975.470 4.280 ;
        RECT 976.310 3.670 978.690 4.280 ;
        RECT 979.530 3.670 982.370 4.280 ;
        RECT 983.210 3.670 985.590 4.280 ;
        RECT 986.430 3.670 989.270 4.280 ;
        RECT 990.110 3.670 992.490 4.280 ;
        RECT 993.330 3.670 995.710 4.280 ;
        RECT 996.550 3.670 999.390 4.280 ;
        RECT 1000.230 3.670 1002.610 4.280 ;
        RECT 1003.450 3.670 1006.290 4.280 ;
        RECT 1007.130 3.670 1009.510 4.280 ;
        RECT 1010.350 3.670 1013.190 4.280 ;
        RECT 1014.030 3.670 1016.410 4.280 ;
        RECT 1017.250 3.670 1020.090 4.280 ;
        RECT 1020.930 3.670 1023.310 4.280 ;
        RECT 1024.150 3.670 1026.990 4.280 ;
        RECT 1027.830 3.670 1030.210 4.280 ;
        RECT 1031.050 3.670 1033.430 4.280 ;
        RECT 1034.270 3.670 1037.110 4.280 ;
        RECT 1037.950 3.670 1040.330 4.280 ;
        RECT 1041.170 3.670 1044.010 4.280 ;
        RECT 1044.850 3.670 1047.230 4.280 ;
        RECT 1048.070 3.670 1050.910 4.280 ;
        RECT 1051.750 3.670 1054.130 4.280 ;
        RECT 1054.970 3.670 1057.810 4.280 ;
        RECT 1058.650 3.670 1061.030 4.280 ;
        RECT 1061.870 3.670 1064.710 4.280 ;
        RECT 1065.550 3.670 1067.930 4.280 ;
        RECT 1068.770 3.670 1071.610 4.280 ;
        RECT 1072.450 3.670 1074.830 4.280 ;
        RECT 1075.670 3.670 1078.050 4.280 ;
        RECT 1078.890 3.670 1081.730 4.280 ;
        RECT 1082.570 3.670 1084.950 4.280 ;
        RECT 1085.790 3.670 1088.630 4.280 ;
        RECT 1089.470 3.670 1091.850 4.280 ;
        RECT 1092.690 3.670 1095.530 4.280 ;
        RECT 1096.370 3.670 1098.750 4.280 ;
        RECT 1099.590 3.670 1102.430 4.280 ;
        RECT 1103.270 3.670 1105.650 4.280 ;
        RECT 1106.490 3.670 1109.330 4.280 ;
        RECT 1110.170 3.670 1112.550 4.280 ;
        RECT 1113.390 3.670 1115.770 4.280 ;
        RECT 1116.610 3.670 1119.450 4.280 ;
        RECT 1120.290 3.670 1122.670 4.280 ;
        RECT 1123.510 3.670 1126.350 4.280 ;
        RECT 1127.190 3.670 1129.570 4.280 ;
        RECT 1130.410 3.670 1133.250 4.280 ;
        RECT 1134.090 3.670 1136.470 4.280 ;
        RECT 1137.310 3.670 1140.150 4.280 ;
        RECT 1140.990 3.670 1143.370 4.280 ;
        RECT 1144.210 3.670 1147.050 4.280 ;
        RECT 1147.890 3.670 1150.270 4.280 ;
        RECT 1151.110 3.670 1153.950 4.280 ;
        RECT 1154.790 3.670 1157.170 4.280 ;
        RECT 1158.010 3.670 1160.390 4.280 ;
        RECT 1161.230 3.670 1164.070 4.280 ;
        RECT 1164.910 3.670 1167.290 4.280 ;
        RECT 1168.130 3.670 1170.970 4.280 ;
        RECT 1171.810 3.670 1174.190 4.280 ;
        RECT 1175.030 3.670 1177.870 4.280 ;
        RECT 1178.710 3.670 1181.090 4.280 ;
        RECT 1181.930 3.670 1184.770 4.280 ;
        RECT 1185.610 3.670 1187.990 4.280 ;
        RECT 1188.830 3.670 1191.670 4.280 ;
        RECT 1192.510 3.670 1194.890 4.280 ;
        RECT 1195.730 3.670 1198.110 4.280 ;
        RECT 1198.950 3.670 1201.790 4.280 ;
        RECT 1202.630 3.670 1205.010 4.280 ;
        RECT 1205.850 3.670 1208.690 4.280 ;
        RECT 1209.530 3.670 1211.910 4.280 ;
        RECT 1212.750 3.670 1215.590 4.280 ;
        RECT 1216.430 3.670 1218.810 4.280 ;
        RECT 1219.650 3.670 1222.490 4.280 ;
        RECT 1223.330 3.670 1225.710 4.280 ;
        RECT 1226.550 3.670 1229.390 4.280 ;
        RECT 1230.230 3.670 1232.610 4.280 ;
        RECT 1233.450 3.670 1236.290 4.280 ;
        RECT 1237.130 3.670 1239.510 4.280 ;
        RECT 1240.350 3.670 1242.730 4.280 ;
        RECT 1243.570 3.670 1246.410 4.280 ;
        RECT 1247.250 3.670 1249.630 4.280 ;
        RECT 1250.470 3.670 1253.310 4.280 ;
        RECT 1254.150 3.670 1256.530 4.280 ;
        RECT 1257.370 3.670 1260.210 4.280 ;
        RECT 1261.050 3.670 1263.430 4.280 ;
        RECT 1264.270 3.670 1267.110 4.280 ;
        RECT 1267.950 3.670 1270.330 4.280 ;
        RECT 1271.170 3.670 1274.010 4.280 ;
        RECT 1274.850 3.670 1277.230 4.280 ;
        RECT 1278.070 3.670 1280.450 4.280 ;
        RECT 1281.290 3.670 1284.130 4.280 ;
        RECT 1284.970 3.670 1287.350 4.280 ;
        RECT 1288.190 3.670 1291.030 4.280 ;
        RECT 1291.870 3.670 1294.250 4.280 ;
        RECT 1295.090 3.670 1297.930 4.280 ;
        RECT 1298.770 3.670 1301.150 4.280 ;
        RECT 1301.990 3.670 1304.830 4.280 ;
        RECT 1305.670 3.670 1308.050 4.280 ;
        RECT 1308.890 3.670 1311.730 4.280 ;
        RECT 1312.570 3.670 1314.950 4.280 ;
        RECT 1315.790 3.670 1318.630 4.280 ;
        RECT 1319.470 3.670 1321.850 4.280 ;
        RECT 1322.690 3.670 1325.070 4.280 ;
        RECT 1325.910 3.670 1328.750 4.280 ;
        RECT 1329.590 3.670 1331.970 4.280 ;
        RECT 1332.810 3.670 1335.650 4.280 ;
        RECT 1336.490 3.670 1338.870 4.280 ;
        RECT 1339.710 3.670 1342.550 4.280 ;
        RECT 1343.390 3.670 1345.770 4.280 ;
        RECT 1346.610 3.670 1349.450 4.280 ;
        RECT 1350.290 3.670 1352.670 4.280 ;
        RECT 1353.510 3.670 1356.350 4.280 ;
        RECT 1357.190 3.670 1359.570 4.280 ;
        RECT 1360.410 3.670 1362.790 4.280 ;
        RECT 1363.630 3.670 1366.470 4.280 ;
        RECT 1367.310 3.670 1369.690 4.280 ;
        RECT 1370.530 3.670 1373.370 4.280 ;
        RECT 1374.210 3.670 1376.590 4.280 ;
        RECT 1377.430 3.670 1380.270 4.280 ;
        RECT 1381.110 3.670 1383.490 4.280 ;
        RECT 1384.330 3.670 1387.170 4.280 ;
        RECT 1388.010 3.670 1390.390 4.280 ;
        RECT 1391.230 3.670 1394.070 4.280 ;
        RECT 1394.910 3.670 1397.290 4.280 ;
        RECT 1398.130 3.670 1400.970 4.280 ;
        RECT 1401.810 3.670 1404.190 4.280 ;
        RECT 1405.030 3.670 1407.410 4.280 ;
        RECT 1408.250 3.670 1411.090 4.280 ;
        RECT 1411.930 3.670 1414.310 4.280 ;
        RECT 1415.150 3.670 1417.990 4.280 ;
        RECT 1418.830 3.670 1421.210 4.280 ;
        RECT 1422.050 3.670 1424.890 4.280 ;
        RECT 1425.730 3.670 1428.110 4.280 ;
        RECT 1428.950 3.670 1431.790 4.280 ;
        RECT 1432.630 3.670 1435.010 4.280 ;
        RECT 1435.850 3.670 1438.690 4.280 ;
        RECT 1439.530 3.670 1441.910 4.280 ;
        RECT 1442.750 3.670 1445.130 4.280 ;
        RECT 1445.970 3.670 1448.810 4.280 ;
        RECT 1449.650 3.670 1452.030 4.280 ;
        RECT 1452.870 3.670 1455.710 4.280 ;
        RECT 1456.550 3.670 1458.930 4.280 ;
        RECT 1459.770 3.670 1462.610 4.280 ;
        RECT 1463.450 3.670 1465.830 4.280 ;
        RECT 1466.670 3.670 1469.510 4.280 ;
        RECT 1470.350 3.670 1472.730 4.280 ;
        RECT 1473.570 3.670 1476.410 4.280 ;
        RECT 1477.250 3.670 1479.630 4.280 ;
        RECT 1480.470 3.670 1483.310 4.280 ;
        RECT 1484.150 3.670 1486.530 4.280 ;
        RECT 1487.370 3.670 1489.750 4.280 ;
        RECT 1490.590 3.670 1493.430 4.280 ;
        RECT 1494.270 3.670 1496.650 4.280 ;
        RECT 1497.490 3.670 1500.330 4.280 ;
        RECT 1501.170 3.670 1503.550 4.280 ;
        RECT 1504.390 3.670 1507.230 4.280 ;
        RECT 1508.070 3.670 1510.450 4.280 ;
        RECT 1511.290 3.670 1514.130 4.280 ;
        RECT 1514.970 3.670 1517.350 4.280 ;
        RECT 1518.190 3.670 1521.030 4.280 ;
        RECT 1521.870 3.670 1524.250 4.280 ;
        RECT 1525.090 3.670 1527.470 4.280 ;
        RECT 1528.310 3.670 1531.150 4.280 ;
        RECT 1531.990 3.670 1534.370 4.280 ;
        RECT 1535.210 3.670 1538.050 4.280 ;
        RECT 1538.890 3.670 1541.270 4.280 ;
        RECT 1542.110 3.670 1544.950 4.280 ;
        RECT 1545.790 3.670 1548.170 4.280 ;
        RECT 1549.010 3.670 1551.850 4.280 ;
        RECT 1552.690 3.670 1555.070 4.280 ;
        RECT 1555.910 3.670 1558.750 4.280 ;
        RECT 1559.590 3.670 1561.970 4.280 ;
        RECT 1562.810 3.670 1565.650 4.280 ;
        RECT 1566.490 3.670 1568.870 4.280 ;
        RECT 1569.710 3.670 1572.090 4.280 ;
        RECT 1572.930 3.670 1575.770 4.280 ;
        RECT 1576.610 3.670 1578.990 4.280 ;
        RECT 1579.830 3.670 1582.670 4.280 ;
        RECT 1583.510 3.670 1585.890 4.280 ;
        RECT 1586.730 3.670 1589.570 4.280 ;
        RECT 1590.410 3.670 1592.790 4.280 ;
        RECT 1593.630 3.670 1596.470 4.280 ;
        RECT 1597.310 3.670 1599.690 4.280 ;
        RECT 1600.530 3.670 1603.370 4.280 ;
        RECT 1604.210 3.670 1606.590 4.280 ;
        RECT 1607.430 3.670 1609.810 4.280 ;
        RECT 1610.650 3.670 1613.490 4.280 ;
        RECT 1614.330 3.670 1616.710 4.280 ;
        RECT 1617.550 3.670 1620.390 4.280 ;
        RECT 1621.230 3.670 1623.610 4.280 ;
        RECT 1624.450 3.670 1627.290 4.280 ;
        RECT 1628.130 3.670 1630.510 4.280 ;
        RECT 1631.350 3.670 1634.190 4.280 ;
        RECT 1635.030 3.670 1637.410 4.280 ;
        RECT 1638.250 3.670 1641.090 4.280 ;
        RECT 1641.930 3.670 1644.310 4.280 ;
        RECT 1645.150 3.670 1647.990 4.280 ;
        RECT 1648.830 3.670 1651.210 4.280 ;
        RECT 1652.050 3.670 1654.430 4.280 ;
        RECT 1655.270 3.670 1658.110 4.280 ;
        RECT 1658.950 3.670 1661.330 4.280 ;
        RECT 1662.170 3.670 1665.010 4.280 ;
        RECT 1665.850 3.670 1668.230 4.280 ;
        RECT 1669.070 3.670 1671.910 4.280 ;
        RECT 1672.750 3.670 1675.130 4.280 ;
        RECT 1675.970 3.670 1678.810 4.280 ;
        RECT 1679.650 3.670 1682.030 4.280 ;
        RECT 1682.870 3.670 1685.710 4.280 ;
        RECT 1686.550 3.670 1688.930 4.280 ;
      LAYER met3 ;
        RECT 21.040 9.015 1656.395 2026.565 ;
      LAYER met4 ;
        RECT 265.255 18.535 327.840 2008.545 ;
        RECT 330.240 18.535 404.640 2008.545 ;
        RECT 407.040 18.535 481.440 2008.545 ;
        RECT 483.840 18.535 558.240 2008.545 ;
        RECT 560.640 18.535 635.040 2008.545 ;
        RECT 637.440 18.535 711.840 2008.545 ;
        RECT 714.240 18.535 788.640 2008.545 ;
        RECT 791.040 18.535 865.440 2008.545 ;
        RECT 867.840 18.535 942.240 2008.545 ;
        RECT 944.640 18.535 1019.040 2008.545 ;
        RECT 1021.440 18.535 1095.840 2008.545 ;
        RECT 1098.240 18.535 1172.640 2008.545 ;
        RECT 1175.040 18.535 1249.440 2008.545 ;
        RECT 1251.840 18.535 1326.240 2008.545 ;
        RECT 1328.640 18.535 1403.040 2008.545 ;
        RECT 1405.440 18.535 1479.840 2008.545 ;
        RECT 1482.240 18.535 1556.345 2008.545 ;
  END
END user_project
END LIBRARY

